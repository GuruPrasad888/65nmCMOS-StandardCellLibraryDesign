module INV(IN, OUT);
input IN;
output OUT;
assign OUT = ~IN;
endmodule

module NAND2(A, B, OUT);
input A, B;
output OUT;
assign OUT = ~(A & B);
endmodule

module NAND3(A, B, C, OUT);
input A, B, C;
output OUT;
assign OUT = ~(A & B & C);
endmodule

module NAND4(A, B, C, D, OUT);
input A, B, C, D;
output OUT;
assign OUT = ~(A & B & C & D);
endmodule

module NOR2(A, B, OUT);
input A, B;
output OUT;
assign OUT = ~(A | B);
endmodule

module NOR3(A, B, C, OUT);
input A, B, C;
output OUT;
assign OUT = ~(A | B | C);
endmodule

module XOR2(A, B, OUT);
input A, B;
output OUT;
assign OUT = (A ^ B);
endmodule

module AOI12(A, B, C, OUT);
input A, B, C;
output OUT;
assign OUT = ~(A | (B & C));
endmodule

module AOI22(A, B, C, D, OUT);
input A, B, C, D;
output OUT;
assign OUT = ~((A & B) | (C & D));
endmodule

module OAI12(A, B, C, OUT);
input A, B, C;
output OUT;
assign OUT = ~(A & (B | C));
endmodule

module OAI22(A, B, C, D, OUT);
input A, B, C, D;
output OUT;
assign OUT = ~((A | B) & (C | D));
endmodule

module DFF( D, CLK, R, Q);
input D, CLK, R;
output Q;
reg Q;
always @(negedge CLK or posedge R)
  if (R == 1'b1)
    Q = 1'b0;
  else
    Q = D;
endmodule




module ALU ( clk, A, B, reset_n, select, F );
  input [31:0] A;
  input [31:0] B;
  input [2:0] select;
  output [31:0] F;
  input clk, reset_n;
  wire   N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23,
         N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51,
         N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N78, N79, N80, N82,
         N83, N85, N86, N87, N88, N90, N91, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229,
         N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240,
         N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251,
         N252, N253, n44, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, \mult_49/A1[0] , \mult_49/A1[1] , \mult_49/A1[2] ,
         \mult_49/A1[3] , \mult_49/A1[4] , \mult_49/A1[5] , \mult_49/A1[6] ,
         \mult_49/A1[7] , \mult_49/A1[8] , \mult_49/A1[9] , \mult_49/A1[10] ,
         \mult_49/A1[11] , \mult_49/A1[12] , \mult_49/A1[13] ,
         \mult_49/A1[14] , \mult_49/A1[15] , \mult_49/A1[16] ,
         \mult_49/A1[17] , \mult_49/A1[18] , \mult_49/A1[19] ,
         \mult_49/A1[20] , \mult_49/A1[21] , \mult_49/A1[22] ,
         \mult_49/A1[23] , \mult_49/A1[24] , \mult_49/A1[25] ,
         \mult_49/A1[26] , \mult_49/A1[27] , \mult_49/A1[28] ,
         \mult_49/A1[29] , \mult_49/ab[0][1] , \mult_49/ab[0][2] ,
         \mult_49/ab[0][3] , \mult_49/ab[0][4] , \mult_49/ab[0][5] ,
         \mult_49/ab[0][6] , \mult_49/ab[0][7] , \mult_49/ab[0][8] ,
         \mult_49/ab[0][9] , \mult_49/ab[0][10] , \mult_49/ab[0][11] ,
         \mult_49/ab[0][12] , \mult_49/ab[0][13] , \mult_49/ab[0][14] ,
         \mult_49/ab[0][15] , \mult_49/ab[0][16] , \mult_49/ab[0][17] ,
         \mult_49/ab[0][18] , \mult_49/ab[0][19] , \mult_49/ab[0][20] ,
         \mult_49/ab[0][21] , \mult_49/ab[0][22] , \mult_49/ab[0][23] ,
         \mult_49/ab[0][24] , \mult_49/ab[0][25] , \mult_49/ab[0][26] ,
         \mult_49/ab[0][27] , \mult_49/ab[0][28] , \mult_49/ab[0][29] ,
         \mult_49/ab[0][30] , \mult_49/ab[0][31] , \mult_49/ab[1][0] ,
         \mult_49/ab[1][1] , \mult_49/ab[1][2] , \mult_49/ab[1][3] ,
         \mult_49/ab[1][4] , \mult_49/ab[1][5] , \mult_49/ab[1][6] ,
         \mult_49/ab[1][7] , \mult_49/ab[1][8] , \mult_49/ab[1][9] ,
         \mult_49/ab[1][10] , \mult_49/ab[1][11] , \mult_49/ab[1][12] ,
         \mult_49/ab[1][13] , \mult_49/ab[1][14] , \mult_49/ab[1][15] ,
         \mult_49/ab[1][16] , \mult_49/ab[1][17] , \mult_49/ab[1][18] ,
         \mult_49/ab[1][19] , \mult_49/ab[1][20] , \mult_49/ab[1][21] ,
         \mult_49/ab[1][22] , \mult_49/ab[1][23] , \mult_49/ab[1][24] ,
         \mult_49/ab[1][25] , \mult_49/ab[1][26] , \mult_49/ab[1][27] ,
         \mult_49/ab[1][28] , \mult_49/ab[1][29] , \mult_49/ab[1][30] ,
         \mult_49/ab[2][0] , \mult_49/ab[2][1] , \mult_49/ab[2][2] ,
         \mult_49/ab[2][3] , \mult_49/ab[2][4] , \mult_49/ab[2][5] ,
         \mult_49/ab[2][6] , \mult_49/ab[2][7] , \mult_49/ab[2][8] ,
         \mult_49/ab[2][9] , \mult_49/ab[2][10] , \mult_49/ab[2][11] ,
         \mult_49/ab[2][12] , \mult_49/ab[2][13] , \mult_49/ab[2][14] ,
         \mult_49/ab[2][15] , \mult_49/ab[2][16] , \mult_49/ab[2][17] ,
         \mult_49/ab[2][18] , \mult_49/ab[2][19] , \mult_49/ab[2][20] ,
         \mult_49/ab[2][21] , \mult_49/ab[2][22] , \mult_49/ab[2][23] ,
         \mult_49/ab[2][24] , \mult_49/ab[2][25] , \mult_49/ab[2][26] ,
         \mult_49/ab[2][27] , \mult_49/ab[2][28] , \mult_49/ab[2][29] ,
         \mult_49/ab[3][0] , \mult_49/ab[3][1] , \mult_49/ab[3][2] ,
         \mult_49/ab[3][3] , \mult_49/ab[3][4] , \mult_49/ab[3][5] ,
         \mult_49/ab[3][6] , \mult_49/ab[3][7] , \mult_49/ab[3][8] ,
         \mult_49/ab[3][9] , \mult_49/ab[3][10] , \mult_49/ab[3][11] ,
         \mult_49/ab[3][12] , \mult_49/ab[3][13] , \mult_49/ab[3][14] ,
         \mult_49/ab[3][15] , \mult_49/ab[3][16] , \mult_49/ab[3][17] ,
         \mult_49/ab[3][18] , \mult_49/ab[3][19] , \mult_49/ab[3][20] ,
         \mult_49/ab[3][21] , \mult_49/ab[3][22] , \mult_49/ab[3][23] ,
         \mult_49/ab[3][24] , \mult_49/ab[3][25] , \mult_49/ab[3][26] ,
         \mult_49/ab[3][27] , \mult_49/ab[3][28] , \mult_49/ab[4][0] ,
         \mult_49/ab[4][1] , \mult_49/ab[4][2] , \mult_49/ab[4][3] ,
         \mult_49/ab[4][4] , \mult_49/ab[4][5] , \mult_49/ab[4][6] ,
         \mult_49/ab[4][7] , \mult_49/ab[4][8] , \mult_49/ab[4][9] ,
         \mult_49/ab[4][10] , \mult_49/ab[4][11] , \mult_49/ab[4][12] ,
         \mult_49/ab[4][13] , \mult_49/ab[4][14] , \mult_49/ab[4][15] ,
         \mult_49/ab[4][16] , \mult_49/ab[4][17] , \mult_49/ab[4][18] ,
         \mult_49/ab[4][19] , \mult_49/ab[4][20] , \mult_49/ab[4][21] ,
         \mult_49/ab[4][22] , \mult_49/ab[4][23] , \mult_49/ab[4][24] ,
         \mult_49/ab[4][25] , \mult_49/ab[4][26] , \mult_49/ab[4][27] ,
         \mult_49/ab[5][0] , \mult_49/ab[5][1] , \mult_49/ab[5][2] ,
         \mult_49/ab[5][3] , \mult_49/ab[5][4] , \mult_49/ab[5][5] ,
         \mult_49/ab[5][6] , \mult_49/ab[5][7] , \mult_49/ab[5][8] ,
         \mult_49/ab[5][9] , \mult_49/ab[5][10] , \mult_49/ab[5][11] ,
         \mult_49/ab[5][12] , \mult_49/ab[5][13] , \mult_49/ab[5][14] ,
         \mult_49/ab[5][15] , \mult_49/ab[5][16] , \mult_49/ab[5][17] ,
         \mult_49/ab[5][18] , \mult_49/ab[5][19] , \mult_49/ab[5][20] ,
         \mult_49/ab[5][21] , \mult_49/ab[5][22] , \mult_49/ab[5][23] ,
         \mult_49/ab[5][24] , \mult_49/ab[5][25] , \mult_49/ab[5][26] ,
         \mult_49/ab[6][0] , \mult_49/ab[6][1] , \mult_49/ab[6][2] ,
         \mult_49/ab[6][3] , \mult_49/ab[6][4] , \mult_49/ab[6][5] ,
         \mult_49/ab[6][6] , \mult_49/ab[6][7] , \mult_49/ab[6][8] ,
         \mult_49/ab[6][9] , \mult_49/ab[6][10] , \mult_49/ab[6][11] ,
         \mult_49/ab[6][12] , \mult_49/ab[6][13] , \mult_49/ab[6][14] ,
         \mult_49/ab[6][15] , \mult_49/ab[6][16] , \mult_49/ab[6][17] ,
         \mult_49/ab[6][18] , \mult_49/ab[6][19] , \mult_49/ab[6][20] ,
         \mult_49/ab[6][21] , \mult_49/ab[6][22] , \mult_49/ab[6][23] ,
         \mult_49/ab[6][24] , \mult_49/ab[6][25] , \mult_49/ab[7][0] ,
         \mult_49/ab[7][1] , \mult_49/ab[7][2] , \mult_49/ab[7][3] ,
         \mult_49/ab[7][4] , \mult_49/ab[7][5] , \mult_49/ab[7][6] ,
         \mult_49/ab[7][7] , \mult_49/ab[7][8] , \mult_49/ab[7][9] ,
         \mult_49/ab[7][10] , \mult_49/ab[7][11] , \mult_49/ab[7][12] ,
         \mult_49/ab[7][13] , \mult_49/ab[7][14] , \mult_49/ab[7][15] ,
         \mult_49/ab[7][16] , \mult_49/ab[7][17] , \mult_49/ab[7][18] ,
         \mult_49/ab[7][19] , \mult_49/ab[7][20] , \mult_49/ab[7][21] ,
         \mult_49/ab[7][22] , \mult_49/ab[7][23] , \mult_49/ab[7][24] ,
         \mult_49/ab[8][0] , \mult_49/ab[8][1] , \mult_49/ab[8][2] ,
         \mult_49/ab[8][3] , \mult_49/ab[8][4] , \mult_49/ab[8][5] ,
         \mult_49/ab[8][6] , \mult_49/ab[8][7] , \mult_49/ab[8][8] ,
         \mult_49/ab[8][9] , \mult_49/ab[8][10] , \mult_49/ab[8][11] ,
         \mult_49/ab[8][12] , \mult_49/ab[8][13] , \mult_49/ab[8][14] ,
         \mult_49/ab[8][15] , \mult_49/ab[8][16] , \mult_49/ab[8][17] ,
         \mult_49/ab[8][18] , \mult_49/ab[8][19] , \mult_49/ab[8][20] ,
         \mult_49/ab[8][21] , \mult_49/ab[8][22] , \mult_49/ab[8][23] ,
         \mult_49/ab[9][0] , \mult_49/ab[9][1] , \mult_49/ab[9][2] ,
         \mult_49/ab[9][3] , \mult_49/ab[9][4] , \mult_49/ab[9][5] ,
         \mult_49/ab[9][6] , \mult_49/ab[9][7] , \mult_49/ab[9][8] ,
         \mult_49/ab[9][9] , \mult_49/ab[9][10] , \mult_49/ab[9][11] ,
         \mult_49/ab[9][12] , \mult_49/ab[9][13] , \mult_49/ab[9][14] ,
         \mult_49/ab[9][15] , \mult_49/ab[9][16] , \mult_49/ab[9][17] ,
         \mult_49/ab[9][18] , \mult_49/ab[9][19] , \mult_49/ab[9][20] ,
         \mult_49/ab[9][21] , \mult_49/ab[9][22] , \mult_49/ab[10][0] ,
         \mult_49/ab[10][1] , \mult_49/ab[10][2] , \mult_49/ab[10][3] ,
         \mult_49/ab[10][4] , \mult_49/ab[10][5] , \mult_49/ab[10][6] ,
         \mult_49/ab[10][7] , \mult_49/ab[10][8] , \mult_49/ab[10][9] ,
         \mult_49/ab[10][10] , \mult_49/ab[10][11] , \mult_49/ab[10][12] ,
         \mult_49/ab[10][13] , \mult_49/ab[10][14] , \mult_49/ab[10][15] ,
         \mult_49/ab[10][16] , \mult_49/ab[10][17] , \mult_49/ab[10][18] ,
         \mult_49/ab[10][19] , \mult_49/ab[10][20] , \mult_49/ab[10][21] ,
         \mult_49/ab[11][0] , \mult_49/ab[11][1] , \mult_49/ab[11][2] ,
         \mult_49/ab[11][3] , \mult_49/ab[11][4] , \mult_49/ab[11][5] ,
         \mult_49/ab[11][6] , \mult_49/ab[11][7] , \mult_49/ab[11][8] ,
         \mult_49/ab[11][9] , \mult_49/ab[11][10] , \mult_49/ab[11][11] ,
         \mult_49/ab[11][12] , \mult_49/ab[11][13] , \mult_49/ab[11][14] ,
         \mult_49/ab[11][15] , \mult_49/ab[11][16] , \mult_49/ab[11][17] ,
         \mult_49/ab[11][18] , \mult_49/ab[11][19] , \mult_49/ab[11][20] ,
         \mult_49/ab[12][0] , \mult_49/ab[12][1] , \mult_49/ab[12][2] ,
         \mult_49/ab[12][3] , \mult_49/ab[12][4] , \mult_49/ab[12][5] ,
         \mult_49/ab[12][6] , \mult_49/ab[12][7] , \mult_49/ab[12][8] ,
         \mult_49/ab[12][9] , \mult_49/ab[12][10] , \mult_49/ab[12][11] ,
         \mult_49/ab[12][12] , \mult_49/ab[12][13] , \mult_49/ab[12][14] ,
         \mult_49/ab[12][15] , \mult_49/ab[12][16] , \mult_49/ab[12][17] ,
         \mult_49/ab[12][18] , \mult_49/ab[12][19] , \mult_49/ab[13][0] ,
         \mult_49/ab[13][1] , \mult_49/ab[13][2] , \mult_49/ab[13][3] ,
         \mult_49/ab[13][4] , \mult_49/ab[13][5] , \mult_49/ab[13][6] ,
         \mult_49/ab[13][7] , \mult_49/ab[13][8] , \mult_49/ab[13][9] ,
         \mult_49/ab[13][10] , \mult_49/ab[13][11] , \mult_49/ab[13][12] ,
         \mult_49/ab[13][13] , \mult_49/ab[13][14] , \mult_49/ab[13][15] ,
         \mult_49/ab[13][16] , \mult_49/ab[13][17] , \mult_49/ab[13][18] ,
         \mult_49/ab[14][0] , \mult_49/ab[14][1] , \mult_49/ab[14][2] ,
         \mult_49/ab[14][3] , \mult_49/ab[14][4] , \mult_49/ab[14][5] ,
         \mult_49/ab[14][6] , \mult_49/ab[14][7] , \mult_49/ab[14][8] ,
         \mult_49/ab[14][9] , \mult_49/ab[14][10] , \mult_49/ab[14][11] ,
         \mult_49/ab[14][12] , \mult_49/ab[14][13] , \mult_49/ab[14][14] ,
         \mult_49/ab[14][15] , \mult_49/ab[14][16] , \mult_49/ab[14][17] ,
         \mult_49/ab[15][0] , \mult_49/ab[15][1] , \mult_49/ab[15][2] ,
         \mult_49/ab[15][3] , \mult_49/ab[15][4] , \mult_49/ab[15][5] ,
         \mult_49/ab[15][6] , \mult_49/ab[15][7] , \mult_49/ab[15][8] ,
         \mult_49/ab[15][9] , \mult_49/ab[15][10] , \mult_49/ab[15][11] ,
         \mult_49/ab[15][12] , \mult_49/ab[15][13] , \mult_49/ab[15][14] ,
         \mult_49/ab[15][15] , \mult_49/ab[15][16] , \mult_49/A_notx[0] ,
         \mult_49/B_notx[0] , \mult_49/ab[16][0] , \mult_49/ab[16][1] ,
         \mult_49/ab[16][2] , \mult_49/ab[16][3] , \mult_49/ab[16][4] ,
         \mult_49/ab[16][5] , \mult_49/ab[16][6] , \mult_49/ab[16][7] ,
         \mult_49/ab[16][8] , \mult_49/ab[16][9] , \mult_49/ab[16][10] ,
         \mult_49/ab[16][11] , \mult_49/ab[16][12] , \mult_49/ab[16][13] ,
         \mult_49/ab[16][14] , \mult_49/ab[16][15] , \mult_49/ab[17][0] ,
         \mult_49/ab[17][1] , \mult_49/ab[17][2] , \mult_49/ab[17][3] ,
         \mult_49/ab[17][4] , \mult_49/ab[17][5] , \mult_49/ab[17][6] ,
         \mult_49/ab[17][7] , \mult_49/ab[17][8] , \mult_49/ab[17][9] ,
         \mult_49/ab[17][10] , \mult_49/ab[17][11] , \mult_49/ab[17][12] ,
         \mult_49/ab[17][13] , \mult_49/ab[17][14] , \mult_49/ab[18][0] ,
         \mult_49/ab[18][1] , \mult_49/ab[18][2] , \mult_49/ab[18][3] ,
         \mult_49/ab[18][4] , \mult_49/ab[18][5] , \mult_49/ab[18][6] ,
         \mult_49/ab[18][7] , \mult_49/ab[18][8] , \mult_49/ab[18][9] ,
         \mult_49/ab[18][10] , \mult_49/ab[18][11] , \mult_49/ab[18][12] ,
         \mult_49/ab[18][13] , \mult_49/ab[19][0] , \mult_49/ab[19][1] ,
         \mult_49/ab[19][2] , \mult_49/ab[19][3] , \mult_49/ab[19][4] ,
         \mult_49/ab[19][5] , \mult_49/ab[19][6] , \mult_49/ab[19][7] ,
         \mult_49/ab[19][8] , \mult_49/ab[19][9] , \mult_49/ab[19][10] ,
         \mult_49/ab[19][11] , \mult_49/ab[19][12] , \mult_49/ab[20][0] ,
         \mult_49/ab[20][1] , \mult_49/ab[20][2] , \mult_49/ab[20][3] ,
         \mult_49/ab[20][4] , \mult_49/ab[20][5] , \mult_49/ab[20][6] ,
         \mult_49/ab[20][7] , \mult_49/ab[20][8] , \mult_49/ab[20][9] ,
         \mult_49/ab[20][10] , \mult_49/ab[20][11] , \mult_49/ab[21][0] ,
         \mult_49/ab[21][1] , \mult_49/ab[21][2] , \mult_49/ab[21][3] ,
         \mult_49/ab[21][4] , \mult_49/ab[21][5] , \mult_49/ab[21][6] ,
         \mult_49/ab[21][7] , \mult_49/ab[21][8] , \mult_49/ab[21][9] ,
         \mult_49/ab[21][10] , \mult_49/ab[22][0] , \mult_49/ab[22][1] ,
         \mult_49/ab[22][2] , \mult_49/ab[22][3] , \mult_49/ab[22][4] ,
         \mult_49/ab[22][5] , \mult_49/ab[22][6] , \mult_49/ab[22][7] ,
         \mult_49/ab[22][8] , \mult_49/ab[22][9] , \mult_49/ab[23][0] ,
         \mult_49/ab[23][1] , \mult_49/ab[23][2] , \mult_49/ab[23][3] ,
         \mult_49/ab[23][4] , \mult_49/ab[23][5] , \mult_49/ab[23][6] ,
         \mult_49/ab[23][7] , \mult_49/ab[23][8] , \mult_49/ab[24][0] ,
         \mult_49/ab[24][1] , \mult_49/ab[24][2] , \mult_49/ab[24][3] ,
         \mult_49/ab[24][4] , \mult_49/ab[24][5] , \mult_49/ab[24][6] ,
         \mult_49/ab[24][7] , \mult_49/ab[25][0] , \mult_49/ab[25][1] ,
         \mult_49/ab[25][2] , \mult_49/ab[25][3] , \mult_49/ab[25][4] ,
         \mult_49/ab[25][5] , \mult_49/ab[25][6] , \mult_49/ab[26][0] ,
         \mult_49/ab[26][1] , \mult_49/ab[26][2] , \mult_49/ab[26][3] ,
         \mult_49/ab[26][4] , \mult_49/ab[26][5] , \mult_49/ab[27][0] ,
         \mult_49/ab[27][1] , \mult_49/ab[27][2] , \mult_49/ab[27][3] ,
         \mult_49/ab[27][4] , \mult_49/ab[28][0] , \mult_49/ab[28][1] ,
         \mult_49/ab[28][2] , \mult_49/ab[28][3] , \mult_49/ab[29][0] ,
         \mult_49/ab[29][1] , \mult_49/ab[29][2] , \mult_49/ab[30][0] ,
         \mult_49/ab[30][1] , \mult_49/ab[31][0] , \gt_48/SB , \gt_48/SA ,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492;
  wire   [31:0] \mult_49/B_not ;
  wire   [31:0] \mult_49/A_not ;
  wire   [31:0] \gt_48/LTV2 ;
  wire   [31:0] \gt_48/LTV1 ;
  wire   [31:0] \gt_48/AEQB ;
  wire   [31:1] \gt_48/LTV ;
  assign \gt_48/SB  = A[31];
  assign \gt_48/SA  = B[31];

  INV I_72 ( .IN(A[0]), .OUT(N220) );
  INV I_40 ( .IN(N90), .OUT(N91) );
  INV I_39 ( .IN(N87), .OUT(N88) );
  INV I_38 ( .IN(N85), .OUT(N86) );
  INV I_36 ( .IN(N82), .OUT(N83) );
  INV I_35 ( .IN(select[1]), .OUT(N80) );
  INV I_34 ( .IN(N78), .OUT(N79) );
  INV I_33 ( .IN(select[2]), .OUT(N74) );
  INV I_32 ( .IN(B[0]), .OUT(N73) );
  INV I_31 ( .IN(B[1]), .OUT(N72) );
  INV I_30 ( .IN(B[2]), .OUT(N71) );
  INV I_29 ( .IN(B[3]), .OUT(N70) );
  INV I_28 ( .IN(B[4]), .OUT(N69) );
  INV I_27 ( .IN(B[5]), .OUT(N68) );
  INV I_26 ( .IN(B[6]), .OUT(N67) );
  INV I_25 ( .IN(B[7]), .OUT(N66) );
  INV I_24 ( .IN(B[8]), .OUT(N65) );
  INV I_23 ( .IN(B[9]), .OUT(N64) );
  INV I_22 ( .IN(B[10]), .OUT(N63) );
  INV I_21 ( .IN(B[11]), .OUT(N62) );
  INV I_20 ( .IN(B[12]), .OUT(N61) );
  INV I_19 ( .IN(B[13]), .OUT(N60) );
  INV I_18 ( .IN(B[14]), .OUT(N59) );
  INV I_17 ( .IN(B[15]), .OUT(N58) );
  INV I_16 ( .IN(B[16]), .OUT(N57) );
  INV I_15 ( .IN(B[17]), .OUT(N56) );
  INV I_14 ( .IN(B[18]), .OUT(N55) );
  INV I_13 ( .IN(B[19]), .OUT(N54) );
  INV I_12 ( .IN(B[20]), .OUT(N53) );
  INV I_11 ( .IN(B[21]), .OUT(N52) );
  INV I_10 ( .IN(B[22]), .OUT(N51) );
  INV I_9 ( .IN(B[23]), .OUT(N50) );
  INV I_8 ( .IN(B[24]), .OUT(N49) );
  INV I_7 ( .IN(B[25]), .OUT(N48) );
  INV I_6 ( .IN(B[26]), .OUT(N47) );
  INV I_5 ( .IN(B[27]), .OUT(N46) );
  INV I_4 ( .IN(B[28]), .OUT(N45) );
  INV I_3 ( .IN(B[29]), .OUT(N44) );
  INV I_2 ( .IN(B[30]), .OUT(N43) );
  INV I_1 ( .IN(\gt_48/SA ), .OUT(N42) );
  NOR2 C97 ( .A(N74), .B(select[1]), .OUT(n46) );
  NOR2 C83 ( .A(select[2]), .B(N80), .OUT(n47) );
  NOR2 C79 ( .A(select[2]), .B(select[1]), .OUT(n48) );
  NOR2 C76 ( .A(select[2]), .B(select[1]), .OUT(N75) );
  DFF \F_out_reg[31]  ( .D(N41), .CLK(n44), .R(1'b0), .Q(F[31]) );
  DFF \F_out_reg[30]  ( .D(N40), .CLK(n44), .R(1'b0), .Q(F[30]) );
  DFF \F_out_reg[29]  ( .D(N39), .CLK(n44), .R(1'b0), .Q(F[29]) );
  DFF \F_out_reg[28]  ( .D(N38), .CLK(n44), .R(1'b0), .Q(F[28]) );
  DFF \F_out_reg[27]  ( .D(N37), .CLK(n44), .R(1'b0), .Q(F[27]) );
  DFF \F_out_reg[26]  ( .D(N36), .CLK(n44), .R(1'b0), .Q(F[26]) );
  DFF \F_out_reg[25]  ( .D(N35), .CLK(n44), .R(1'b0), .Q(F[25]) );
  DFF \F_out_reg[24]  ( .D(N34), .CLK(n44), .R(1'b0), .Q(F[24]) );
  DFF \F_out_reg[23]  ( .D(N33), .CLK(n44), .R(1'b0), .Q(F[23]) );
  DFF \F_out_reg[22]  ( .D(N32), .CLK(n44), .R(1'b0), .Q(F[22]) );
  DFF \F_out_reg[21]  ( .D(N31), .CLK(n44), .R(1'b0), .Q(F[21]) );
  DFF \F_out_reg[20]  ( .D(N30), .CLK(n44), .R(1'b0), .Q(F[20]) );
  DFF \F_out_reg[19]  ( .D(N29), .CLK(n44), .R(1'b0), .Q(F[19]) );
  DFF \F_out_reg[18]  ( .D(N28), .CLK(n44), .R(1'b0), .Q(F[18]) );
  DFF \F_out_reg[17]  ( .D(N27), .CLK(n44), .R(1'b0), .Q(F[17]) );
  DFF \F_out_reg[16]  ( .D(N26), .CLK(n44), .R(1'b0), .Q(F[16]) );
  DFF \F_out_reg[15]  ( .D(N25), .CLK(n44), .R(1'b0), .Q(F[15]) );
  DFF \F_out_reg[14]  ( .D(N24), .CLK(n44), .R(1'b0), .Q(F[14]) );
  DFF \F_out_reg[13]  ( .D(N23), .CLK(n44), .R(1'b0), .Q(F[13]) );
  DFF \F_out_reg[12]  ( .D(N22), .CLK(n44), .R(1'b0), .Q(F[12]) );
  DFF \F_out_reg[11]  ( .D(N21), .CLK(n44), .R(1'b0), .Q(F[11]) );
  DFF \F_out_reg[10]  ( .D(N20), .CLK(n44), .R(1'b0), .Q(F[10]) );
  DFF \F_out_reg[9]  ( .D(N19), .CLK(n44), .R(1'b0), .Q(F[9]) );
  DFF \F_out_reg[8]  ( .D(N18), .CLK(n44), .R(1'b0), .Q(F[8]) );
  DFF \F_out_reg[7]  ( .D(N17), .CLK(n44), .R(1'b0), .Q(F[7]) );
  DFF \F_out_reg[6]  ( .D(N16), .CLK(n44), .R(1'b0), .Q(F[6]) );
  DFF \F_out_reg[5]  ( .D(N15), .CLK(n44), .R(1'b0), .Q(F[5]) );
  DFF \F_out_reg[4]  ( .D(N14), .CLK(n44), .R(1'b0), .Q(F[4]) );
  DFF \F_out_reg[3]  ( .D(N13), .CLK(n44), .R(1'b0), .Q(F[3]) );
  DFF \F_out_reg[2]  ( .D(N12), .CLK(n44), .R(1'b0), .Q(F[2]) );
  DFF \F_out_reg[1]  ( .D(N11), .CLK(n44), .R(1'b0), .Q(F[1]) );
  DFF \F_out_reg[0]  ( .D(N10), .CLK(n44), .R(1'b0), .Q(F[0]) );
  INV U37 ( .IN(clk), .OUT(n44) );
  NAND2 U39 ( .A(select[0]), .B(n46), .OUT(N90) );
  NAND2 U40 ( .A(n46), .B(n49), .OUT(N87) );
  NAND2 U41 ( .A(n47), .B(select[0]), .OUT(N85) );
  NAND2 U42 ( .A(n47), .B(n49), .OUT(N82) );
  NAND2 U43 ( .A(n48), .B(select[0]), .OUT(N78) );
  NAND3 U44 ( .A(n50), .B(n51), .C(n52), .OUT(N41) );
  NOR2 U45 ( .A(n53), .B(n54), .OUT(n52) );
  NAND2 U46 ( .A(n55), .B(n56), .OUT(n54) );
  NAND2 U47 ( .A(N124), .B(n57), .OUT(n56) );
  NAND2 U48 ( .A(N188), .B(n58), .OUT(n55) );
  NOR2 U49 ( .A(n59), .B(\gt_48/SB ), .OUT(n53) );
  NAND2 U50 ( .A(N42), .B(n60), .OUT(n51) );
  NAND2 U51 ( .A(N253), .B(n61), .OUT(n50) );
  NAND3 U52 ( .A(n62), .B(n63), .C(n64), .OUT(N40) );
  NOR2 U53 ( .A(n65), .B(n66), .OUT(n64) );
  NAND2 U54 ( .A(n67), .B(n68), .OUT(n66) );
  NAND2 U55 ( .A(N123), .B(n57), .OUT(n68) );
  NAND2 U56 ( .A(N187), .B(n58), .OUT(n67) );
  NOR2 U57 ( .A(n59), .B(A[30]), .OUT(n65) );
  NAND2 U58 ( .A(N43), .B(n60), .OUT(n63) );
  NAND2 U59 ( .A(N252), .B(n61), .OUT(n62) );
  NAND3 U60 ( .A(n69), .B(n70), .C(n71), .OUT(N39) );
  NOR2 U61 ( .A(n72), .B(n73), .OUT(n71) );
  NAND2 U62 ( .A(n74), .B(n75), .OUT(n73) );
  NAND2 U63 ( .A(N122), .B(n57), .OUT(n75) );
  NAND2 U64 ( .A(N186), .B(n58), .OUT(n74) );
  NOR2 U65 ( .A(n59), .B(A[29]), .OUT(n72) );
  NAND2 U66 ( .A(N44), .B(n60), .OUT(n70) );
  NAND2 U67 ( .A(N251), .B(n61), .OUT(n69) );
  NAND3 U68 ( .A(n76), .B(n77), .C(n78), .OUT(N38) );
  NOR2 U69 ( .A(n79), .B(n80), .OUT(n78) );
  NAND2 U70 ( .A(n81), .B(n82), .OUT(n80) );
  NAND2 U71 ( .A(N121), .B(n57), .OUT(n82) );
  NAND2 U72 ( .A(N185), .B(n58), .OUT(n81) );
  NOR2 U73 ( .A(n59), .B(A[28]), .OUT(n79) );
  NAND2 U74 ( .A(N45), .B(n60), .OUT(n77) );
  NAND2 U75 ( .A(N250), .B(n61), .OUT(n76) );
  NAND3 U76 ( .A(n83), .B(n84), .C(n85), .OUT(N37) );
  NOR2 U77 ( .A(n86), .B(n87), .OUT(n85) );
  NAND2 U78 ( .A(n88), .B(n89), .OUT(n87) );
  NAND2 U79 ( .A(N120), .B(n57), .OUT(n89) );
  NAND2 U80 ( .A(N184), .B(n58), .OUT(n88) );
  NOR2 U81 ( .A(n59), .B(A[27]), .OUT(n86) );
  NAND2 U82 ( .A(N46), .B(n60), .OUT(n84) );
  NAND2 U83 ( .A(N249), .B(n61), .OUT(n83) );
  NAND3 U84 ( .A(n90), .B(n91), .C(n92), .OUT(N36) );
  NOR2 U85 ( .A(n93), .B(n94), .OUT(n92) );
  NAND2 U86 ( .A(n95), .B(n96), .OUT(n94) );
  NAND2 U87 ( .A(N119), .B(n57), .OUT(n96) );
  NAND2 U88 ( .A(N183), .B(n58), .OUT(n95) );
  NOR2 U89 ( .A(n59), .B(A[26]), .OUT(n93) );
  NAND2 U90 ( .A(N47), .B(n60), .OUT(n91) );
  NAND2 U91 ( .A(N248), .B(n61), .OUT(n90) );
  NAND3 U92 ( .A(n97), .B(n98), .C(n99), .OUT(N35) );
  NOR2 U93 ( .A(n100), .B(n101), .OUT(n99) );
  NAND2 U94 ( .A(n102), .B(n103), .OUT(n101) );
  NAND2 U95 ( .A(N118), .B(n57), .OUT(n103) );
  NAND2 U96 ( .A(N182), .B(n58), .OUT(n102) );
  NOR2 U97 ( .A(n59), .B(A[25]), .OUT(n100) );
  NAND2 U98 ( .A(N48), .B(n60), .OUT(n98) );
  NAND2 U99 ( .A(N247), .B(n61), .OUT(n97) );
  NAND3 U100 ( .A(n104), .B(n105), .C(n106), .OUT(N34) );
  NOR2 U101 ( .A(n107), .B(n108), .OUT(n106) );
  NAND2 U102 ( .A(n109), .B(n110), .OUT(n108) );
  NAND2 U103 ( .A(N117), .B(n57), .OUT(n110) );
  NAND2 U104 ( .A(N181), .B(n58), .OUT(n109) );
  NOR2 U105 ( .A(n59), .B(A[24]), .OUT(n107) );
  NAND2 U106 ( .A(N49), .B(n60), .OUT(n105) );
  NAND2 U107 ( .A(N246), .B(n61), .OUT(n104) );
  NAND3 U108 ( .A(n111), .B(n112), .C(n113), .OUT(N33) );
  NOR2 U109 ( .A(n114), .B(n115), .OUT(n113) );
  NAND2 U110 ( .A(n116), .B(n117), .OUT(n115) );
  NAND2 U111 ( .A(N116), .B(n57), .OUT(n117) );
  NAND2 U112 ( .A(N180), .B(n58), .OUT(n116) );
  NOR2 U113 ( .A(n59), .B(A[23]), .OUT(n114) );
  NAND2 U114 ( .A(N50), .B(n60), .OUT(n112) );
  NAND2 U115 ( .A(N245), .B(n61), .OUT(n111) );
  NAND3 U116 ( .A(n118), .B(n119), .C(n120), .OUT(N32) );
  NOR2 U117 ( .A(n121), .B(n122), .OUT(n120) );
  NAND2 U118 ( .A(n123), .B(n124), .OUT(n122) );
  NAND2 U119 ( .A(N115), .B(n57), .OUT(n124) );
  NAND2 U120 ( .A(N179), .B(n58), .OUT(n123) );
  NOR2 U121 ( .A(n59), .B(A[22]), .OUT(n121) );
  NAND2 U122 ( .A(N51), .B(n60), .OUT(n119) );
  NAND2 U123 ( .A(N244), .B(n61), .OUT(n118) );
  NAND3 U124 ( .A(n125), .B(n126), .C(n127), .OUT(N31) );
  NOR2 U125 ( .A(n128), .B(n129), .OUT(n127) );
  NAND2 U126 ( .A(n130), .B(n131), .OUT(n129) );
  NAND2 U127 ( .A(N114), .B(n57), .OUT(n131) );
  NAND2 U128 ( .A(N178), .B(n58), .OUT(n130) );
  NOR2 U129 ( .A(n59), .B(A[21]), .OUT(n128) );
  NAND2 U130 ( .A(N52), .B(n60), .OUT(n126) );
  NAND2 U131 ( .A(N243), .B(n61), .OUT(n125) );
  NAND3 U132 ( .A(n132), .B(n133), .C(n134), .OUT(N30) );
  NOR2 U133 ( .A(n135), .B(n136), .OUT(n134) );
  NAND2 U134 ( .A(n137), .B(n138), .OUT(n136) );
  NAND2 U135 ( .A(N113), .B(n57), .OUT(n138) );
  NAND2 U136 ( .A(N177), .B(n58), .OUT(n137) );
  NOR2 U137 ( .A(n59), .B(A[20]), .OUT(n135) );
  NAND2 U138 ( .A(N53), .B(n60), .OUT(n133) );
  NAND2 U139 ( .A(N242), .B(n61), .OUT(n132) );
  NAND3 U140 ( .A(n139), .B(n140), .C(n141), .OUT(N29) );
  NOR2 U141 ( .A(n142), .B(n143), .OUT(n141) );
  NAND2 U142 ( .A(n144), .B(n145), .OUT(n143) );
  NAND2 U143 ( .A(N112), .B(n57), .OUT(n145) );
  NAND2 U144 ( .A(N176), .B(n58), .OUT(n144) );
  NOR2 U145 ( .A(n59), .B(A[19]), .OUT(n142) );
  NAND2 U146 ( .A(N54), .B(n60), .OUT(n140) );
  NAND2 U147 ( .A(N241), .B(n61), .OUT(n139) );
  NAND3 U148 ( .A(n146), .B(n147), .C(n148), .OUT(N28) );
  NOR2 U149 ( .A(n149), .B(n150), .OUT(n148) );
  NAND2 U150 ( .A(n151), .B(n152), .OUT(n150) );
  NAND2 U151 ( .A(N111), .B(n57), .OUT(n152) );
  NAND2 U152 ( .A(N175), .B(n58), .OUT(n151) );
  NOR2 U153 ( .A(n59), .B(A[18]), .OUT(n149) );
  NAND2 U154 ( .A(N55), .B(n60), .OUT(n147) );
  NAND2 U155 ( .A(N240), .B(n61), .OUT(n146) );
  NAND3 U156 ( .A(n153), .B(n154), .C(n155), .OUT(N27) );
  NOR2 U157 ( .A(n156), .B(n157), .OUT(n155) );
  NAND2 U158 ( .A(n158), .B(n159), .OUT(n157) );
  NAND2 U159 ( .A(N110), .B(n57), .OUT(n159) );
  NAND2 U160 ( .A(N174), .B(n58), .OUT(n158) );
  NOR2 U161 ( .A(n59), .B(A[17]), .OUT(n156) );
  NAND2 U162 ( .A(N56), .B(n60), .OUT(n154) );
  NAND2 U163 ( .A(N239), .B(n61), .OUT(n153) );
  NAND3 U164 ( .A(n160), .B(n161), .C(n162), .OUT(N26) );
  NOR2 U165 ( .A(n163), .B(n164), .OUT(n162) );
  NAND2 U166 ( .A(n165), .B(n166), .OUT(n164) );
  NAND2 U167 ( .A(N109), .B(n57), .OUT(n166) );
  NAND2 U168 ( .A(N173), .B(n58), .OUT(n165) );
  NOR2 U169 ( .A(n59), .B(A[16]), .OUT(n163) );
  NAND2 U170 ( .A(N57), .B(n60), .OUT(n161) );
  NAND2 U171 ( .A(N238), .B(n61), .OUT(n160) );
  NAND3 U172 ( .A(n167), .B(n168), .C(n169), .OUT(N25) );
  NOR2 U173 ( .A(n170), .B(n171), .OUT(n169) );
  NAND2 U174 ( .A(n172), .B(n173), .OUT(n171) );
  NAND2 U175 ( .A(N108), .B(n57), .OUT(n173) );
  NAND2 U176 ( .A(N172), .B(n58), .OUT(n172) );
  NOR2 U177 ( .A(n59), .B(A[15]), .OUT(n170) );
  NAND2 U178 ( .A(N58), .B(n60), .OUT(n168) );
  NAND2 U179 ( .A(N237), .B(n61), .OUT(n167) );
  NAND3 U180 ( .A(n174), .B(n175), .C(n176), .OUT(N24) );
  NOR2 U181 ( .A(n177), .B(n178), .OUT(n176) );
  NAND2 U182 ( .A(n179), .B(n180), .OUT(n178) );
  NAND2 U183 ( .A(N107), .B(n57), .OUT(n180) );
  NAND2 U184 ( .A(N171), .B(n58), .OUT(n179) );
  NOR2 U185 ( .A(n59), .B(A[14]), .OUT(n177) );
  NAND2 U186 ( .A(N59), .B(n60), .OUT(n175) );
  NAND2 U187 ( .A(N236), .B(n61), .OUT(n174) );
  NAND3 U188 ( .A(n181), .B(n182), .C(n183), .OUT(N23) );
  NOR2 U189 ( .A(n184), .B(n185), .OUT(n183) );
  NAND2 U190 ( .A(n186), .B(n187), .OUT(n185) );
  NAND2 U191 ( .A(N106), .B(n57), .OUT(n187) );
  NAND2 U192 ( .A(N170), .B(n58), .OUT(n186) );
  NOR2 U193 ( .A(n59), .B(A[13]), .OUT(n184) );
  NAND2 U194 ( .A(N60), .B(n60), .OUT(n182) );
  NAND2 U195 ( .A(N235), .B(n61), .OUT(n181) );
  NAND3 U196 ( .A(n188), .B(n189), .C(n190), .OUT(N22) );
  NOR2 U197 ( .A(n191), .B(n192), .OUT(n190) );
  NAND2 U198 ( .A(n193), .B(n194), .OUT(n192) );
  NAND2 U199 ( .A(N105), .B(n57), .OUT(n194) );
  NAND2 U200 ( .A(N169), .B(n58), .OUT(n193) );
  NOR2 U201 ( .A(n59), .B(A[12]), .OUT(n191) );
  NAND2 U202 ( .A(N61), .B(n60), .OUT(n189) );
  NAND2 U203 ( .A(N234), .B(n61), .OUT(n188) );
  NAND3 U204 ( .A(n195), .B(n196), .C(n197), .OUT(N21) );
  NOR2 U205 ( .A(n198), .B(n199), .OUT(n197) );
  NAND2 U206 ( .A(n200), .B(n201), .OUT(n199) );
  NAND2 U207 ( .A(N104), .B(n57), .OUT(n201) );
  NAND2 U208 ( .A(N168), .B(n58), .OUT(n200) );
  NOR2 U209 ( .A(n59), .B(A[11]), .OUT(n198) );
  NAND2 U210 ( .A(N62), .B(n60), .OUT(n196) );
  NAND2 U211 ( .A(N233), .B(n61), .OUT(n195) );
  NAND3 U212 ( .A(n202), .B(n203), .C(n204), .OUT(N20) );
  NOR2 U213 ( .A(n205), .B(n206), .OUT(n204) );
  NAND2 U214 ( .A(n207), .B(n208), .OUT(n206) );
  NAND2 U215 ( .A(N103), .B(n57), .OUT(n208) );
  NAND2 U216 ( .A(N167), .B(n58), .OUT(n207) );
  NOR2 U217 ( .A(n59), .B(A[10]), .OUT(n205) );
  NAND2 U218 ( .A(N63), .B(n60), .OUT(n203) );
  NAND2 U219 ( .A(N232), .B(n61), .OUT(n202) );
  NAND3 U220 ( .A(n209), .B(n210), .C(n211), .OUT(N19) );
  NOR2 U221 ( .A(n212), .B(n213), .OUT(n211) );
  NAND2 U222 ( .A(n214), .B(n215), .OUT(n213) );
  NAND2 U223 ( .A(N102), .B(n57), .OUT(n215) );
  NAND2 U224 ( .A(N166), .B(n58), .OUT(n214) );
  NOR2 U225 ( .A(n59), .B(A[9]), .OUT(n212) );
  NAND2 U226 ( .A(N64), .B(n60), .OUT(n210) );
  NAND2 U227 ( .A(N231), .B(n61), .OUT(n209) );
  NAND3 U228 ( .A(n216), .B(n217), .C(n218), .OUT(N18) );
  NOR2 U229 ( .A(n219), .B(n220), .OUT(n218) );
  NAND2 U230 ( .A(n221), .B(n222), .OUT(n220) );
  NAND2 U231 ( .A(N101), .B(n57), .OUT(n222) );
  NAND2 U232 ( .A(N165), .B(n58), .OUT(n221) );
  NOR2 U233 ( .A(n59), .B(A[8]), .OUT(n219) );
  NAND2 U234 ( .A(N65), .B(n60), .OUT(n217) );
  NAND2 U235 ( .A(N230), .B(n61), .OUT(n216) );
  NAND3 U236 ( .A(n223), .B(n224), .C(n225), .OUT(N17) );
  NOR2 U237 ( .A(n226), .B(n227), .OUT(n225) );
  NAND2 U238 ( .A(n228), .B(n229), .OUT(n227) );
  NAND2 U239 ( .A(N100), .B(n57), .OUT(n229) );
  NAND2 U240 ( .A(N164), .B(n58), .OUT(n228) );
  NOR2 U241 ( .A(n59), .B(A[7]), .OUT(n226) );
  NAND2 U242 ( .A(N66), .B(n60), .OUT(n224) );
  NAND2 U243 ( .A(N229), .B(n61), .OUT(n223) );
  NAND3 U244 ( .A(n230), .B(n231), .C(n232), .OUT(N16) );
  NOR2 U245 ( .A(n233), .B(n234), .OUT(n232) );
  NAND2 U246 ( .A(n235), .B(n236), .OUT(n234) );
  NAND2 U247 ( .A(N99), .B(n57), .OUT(n236) );
  NAND2 U248 ( .A(N163), .B(n58), .OUT(n235) );
  NOR2 U249 ( .A(n59), .B(A[6]), .OUT(n233) );
  NAND2 U250 ( .A(N67), .B(n60), .OUT(n231) );
  NAND2 U251 ( .A(N228), .B(n61), .OUT(n230) );
  NAND3 U252 ( .A(n237), .B(n238), .C(n239), .OUT(N15) );
  NOR2 U253 ( .A(n240), .B(n241), .OUT(n239) );
  NAND2 U254 ( .A(n242), .B(n243), .OUT(n241) );
  NAND2 U255 ( .A(N98), .B(n57), .OUT(n243) );
  NAND2 U256 ( .A(N162), .B(n58), .OUT(n242) );
  NOR2 U257 ( .A(n59), .B(A[5]), .OUT(n240) );
  NAND2 U258 ( .A(N68), .B(n60), .OUT(n238) );
  NAND2 U259 ( .A(N227), .B(n61), .OUT(n237) );
  NAND3 U260 ( .A(n244), .B(n245), .C(n246), .OUT(N14) );
  NOR2 U261 ( .A(n247), .B(n248), .OUT(n246) );
  NAND2 U262 ( .A(n249), .B(n250), .OUT(n248) );
  NAND2 U263 ( .A(N97), .B(n57), .OUT(n250) );
  NAND2 U264 ( .A(N161), .B(n58), .OUT(n249) );
  NOR2 U265 ( .A(n59), .B(A[4]), .OUT(n247) );
  NAND2 U266 ( .A(N69), .B(n60), .OUT(n245) );
  NAND2 U267 ( .A(N226), .B(n61), .OUT(n244) );
  NAND3 U268 ( .A(n251), .B(n252), .C(n253), .OUT(N13) );
  NOR2 U269 ( .A(n254), .B(n255), .OUT(n253) );
  NAND2 U270 ( .A(n256), .B(n257), .OUT(n255) );
  NAND2 U271 ( .A(N96), .B(n57), .OUT(n257) );
  NAND2 U272 ( .A(N160), .B(n58), .OUT(n256) );
  NOR2 U273 ( .A(n59), .B(A[3]), .OUT(n254) );
  NAND2 U274 ( .A(N70), .B(n60), .OUT(n252) );
  NAND2 U275 ( .A(N225), .B(n61), .OUT(n251) );
  NAND3 U276 ( .A(n258), .B(n259), .C(n260), .OUT(N12) );
  NOR2 U277 ( .A(n261), .B(n262), .OUT(n260) );
  NAND2 U278 ( .A(n263), .B(n264), .OUT(n262) );
  NAND2 U279 ( .A(N95), .B(n57), .OUT(n264) );
  NAND2 U280 ( .A(N159), .B(n58), .OUT(n263) );
  NOR2 U281 ( .A(n59), .B(A[2]), .OUT(n261) );
  NAND2 U282 ( .A(N71), .B(n60), .OUT(n259) );
  NAND2 U283 ( .A(N224), .B(n61), .OUT(n258) );
  NAND3 U284 ( .A(n265), .B(n266), .C(n267), .OUT(N11) );
  NOR2 U285 ( .A(n268), .B(n269), .OUT(n267) );
  NAND2 U286 ( .A(n270), .B(n271), .OUT(n269) );
  NAND2 U287 ( .A(N94), .B(n57), .OUT(n271) );
  NAND2 U288 ( .A(N158), .B(n58), .OUT(n270) );
  NOR2 U289 ( .A(n59), .B(A[1]), .OUT(n268) );
  NAND2 U290 ( .A(N72), .B(n60), .OUT(n266) );
  NAND2 U291 ( .A(N223), .B(n61), .OUT(n265) );
  INV U292 ( .IN(n272), .OUT(N10) );
  NOR2 U293 ( .A(n273), .B(n274), .OUT(n272) );
  NAND3 U294 ( .A(n275), .B(n276), .C(n277), .OUT(n274) );
  NAND2 U295 ( .A(N222), .B(n61), .OUT(n277) );
  INV U296 ( .IN(n278), .OUT(n61) );
  NAND2 U297 ( .A(N91), .B(reset_n), .OUT(n278) );
  NAND2 U298 ( .A(N220), .B(n279), .OUT(n276) );
  INV U299 ( .IN(n59), .OUT(n279) );
  NAND2 U300 ( .A(N83), .B(reset_n), .OUT(n59) );
  NAND2 U301 ( .A(N73), .B(n60), .OUT(n275) );
  INV U302 ( .IN(n280), .OUT(n60) );
  NAND2 U303 ( .A(N86), .B(reset_n), .OUT(n280) );
  NAND3 U304 ( .A(n281), .B(n282), .C(n283), .OUT(n273) );
  NAND2 U305 ( .A(N93), .B(n58), .OUT(n283) );
  INV U306 ( .IN(n284), .OUT(n58) );
  NAND2 U307 ( .A(N79), .B(reset_n), .OUT(n284) );
  NAND3 U308 ( .A(N221), .B(reset_n), .C(N88), .OUT(n282) );
  NAND2 U309 ( .A(N93), .B(n57), .OUT(n281) );
  INV U310 ( .IN(n285), .OUT(n57) );
  NAND2 U311 ( .A(reset_n), .B(n286), .OUT(n285) );
  NAND2 U312 ( .A(n287), .B(n288), .OUT(n286) );
  NAND2 U313 ( .A(N75), .B(n49), .OUT(n288) );
  INV U314 ( .IN(select[0]), .OUT(n49) );
  NAND2 U315 ( .A(select[2]), .B(select[1]), .OUT(n287) );
  INV \mult_49/AN1_31  ( .IN(\gt_48/SB ), .OUT(\mult_49/A_not [31]) );
  INV \mult_49/AN1_30  ( .IN(A[30]), .OUT(\mult_49/A_not [30]) );
  INV \mult_49/AN1_29  ( .IN(A[29]), .OUT(\mult_49/A_not [29]) );
  INV \mult_49/AN1_28  ( .IN(A[28]), .OUT(\mult_49/A_not [28]) );
  INV \mult_49/AN1_27  ( .IN(A[27]), .OUT(\mult_49/A_not [27]) );
  INV \mult_49/AN1_26  ( .IN(A[26]), .OUT(\mult_49/A_not [26]) );
  INV \mult_49/AN1_25  ( .IN(A[25]), .OUT(\mult_49/A_not [25]) );
  INV \mult_49/AN1_24  ( .IN(A[24]), .OUT(\mult_49/A_not [24]) );
  INV \mult_49/AN1_23  ( .IN(A[23]), .OUT(\mult_49/A_not [23]) );
  INV \mult_49/AN1_22  ( .IN(A[22]), .OUT(\mult_49/A_not [22]) );
  INV \mult_49/AN1_21  ( .IN(A[21]), .OUT(\mult_49/A_not [21]) );
  INV \mult_49/AN1_20  ( .IN(A[20]), .OUT(\mult_49/A_not [20]) );
  INV \mult_49/AN1_19  ( .IN(A[19]), .OUT(\mult_49/A_not [19]) );
  INV \mult_49/AN1_18  ( .IN(A[18]), .OUT(\mult_49/A_not [18]) );
  INV \mult_49/AN1_17  ( .IN(A[17]), .OUT(\mult_49/A_not [17]) );
  INV \mult_49/AN1_16  ( .IN(A[16]), .OUT(\mult_49/A_not [16]) );
  INV \mult_49/AN1_15  ( .IN(A[15]), .OUT(\mult_49/A_not [15]) );
  INV \mult_49/AN1_14  ( .IN(A[14]), .OUT(\mult_49/A_not [14]) );
  INV \mult_49/AN1_13  ( .IN(A[13]), .OUT(\mult_49/A_not [13]) );
  INV \mult_49/AN1_12  ( .IN(A[12]), .OUT(\mult_49/A_not [12]) );
  INV \mult_49/AN1_11  ( .IN(A[11]), .OUT(\mult_49/A_not [11]) );
  INV \mult_49/AN1_10  ( .IN(A[10]), .OUT(\mult_49/A_not [10]) );
  INV \mult_49/AN1_9  ( .IN(A[9]), .OUT(\mult_49/A_not [9]) );
  INV \mult_49/AN1_8  ( .IN(A[8]), .OUT(\mult_49/A_not [8]) );
  INV \mult_49/AN1_7  ( .IN(A[7]), .OUT(\mult_49/A_not [7]) );
  INV \mult_49/AN1_6  ( .IN(A[6]), .OUT(\mult_49/A_not [6]) );
  INV \mult_49/AN1_5  ( .IN(A[5]), .OUT(\mult_49/A_not [5]) );
  INV \mult_49/AN1_4  ( .IN(A[4]), .OUT(\mult_49/A_not [4]) );
  INV \mult_49/AN1_3  ( .IN(A[3]), .OUT(\mult_49/A_not [3]) );
  INV \mult_49/AN1_2  ( .IN(A[2]), .OUT(\mult_49/A_not [2]) );
  INV \mult_49/AN1_1  ( .IN(A[1]), .OUT(\mult_49/A_not [1]) );
  INV \mult_49/AN1_0  ( .IN(A[0]), .OUT(\mult_49/A_not [0]) );
  INV \mult_49/AN1_31_0  ( .IN(\gt_48/SA ), .OUT(\mult_49/B_not [31]) );
  INV \mult_49/AN1_30_0  ( .IN(B[30]), .OUT(\mult_49/B_not [30]) );
  INV \mult_49/AN1_29_0  ( .IN(B[29]), .OUT(\mult_49/B_not [29]) );
  INV \mult_49/AN1_28_0  ( .IN(B[28]), .OUT(\mult_49/B_not [28]) );
  INV \mult_49/AN1_27_0  ( .IN(B[27]), .OUT(\mult_49/B_not [27]) );
  INV \mult_49/AN1_26_0  ( .IN(B[26]), .OUT(\mult_49/B_not [26]) );
  INV \mult_49/AN1_25_0  ( .IN(B[25]), .OUT(\mult_49/B_not [25]) );
  INV \mult_49/AN1_24_0  ( .IN(B[24]), .OUT(\mult_49/B_not [24]) );
  INV \mult_49/AN1_23_0  ( .IN(B[23]), .OUT(\mult_49/B_not [23]) );
  INV \mult_49/AN1_22_0  ( .IN(B[22]), .OUT(\mult_49/B_not [22]) );
  INV \mult_49/AN1_21_0  ( .IN(B[21]), .OUT(\mult_49/B_not [21]) );
  INV \mult_49/AN1_20_0  ( .IN(B[20]), .OUT(\mult_49/B_not [20]) );
  INV \mult_49/AN1_19_0  ( .IN(B[19]), .OUT(\mult_49/B_not [19]) );
  INV \mult_49/AN1_18_0  ( .IN(B[18]), .OUT(\mult_49/B_not [18]) );
  INV \mult_49/AN1_17_0  ( .IN(B[17]), .OUT(\mult_49/B_not [17]) );
  INV \mult_49/AN1_16_0  ( .IN(B[16]), .OUT(\mult_49/B_not [16]) );
  INV \mult_49/AN1_15_0  ( .IN(B[15]), .OUT(\mult_49/B_not [15]) );
  INV \mult_49/AN1_14_0  ( .IN(B[14]), .OUT(\mult_49/B_not [14]) );
  INV \mult_49/AN1_13_0  ( .IN(B[13]), .OUT(\mult_49/B_not [13]) );
  INV \mult_49/AN1_12_0  ( .IN(B[12]), .OUT(\mult_49/B_not [12]) );
  INV \mult_49/AN1_11_0  ( .IN(B[11]), .OUT(\mult_49/B_not [11]) );
  INV \mult_49/AN1_10_0  ( .IN(B[10]), .OUT(\mult_49/B_not [10]) );
  INV \mult_49/AN1_9_0  ( .IN(B[9]), .OUT(\mult_49/B_not [9]) );
  INV \mult_49/AN1_8_0  ( .IN(B[8]), .OUT(\mult_49/B_not [8]) );
  INV \mult_49/AN1_7_0  ( .IN(B[7]), .OUT(\mult_49/B_not [7]) );
  INV \mult_49/AN1_6_0  ( .IN(B[6]), .OUT(\mult_49/B_not [6]) );
  INV \mult_49/AN1_5_0  ( .IN(B[5]), .OUT(\mult_49/B_not [5]) );
  INV \mult_49/AN1_4_0  ( .IN(B[4]), .OUT(\mult_49/B_not [4]) );
  INV \mult_49/AN1_3_0  ( .IN(B[3]), .OUT(\mult_49/B_not [3]) );
  INV \mult_49/AN1_2_0  ( .IN(B[2]), .OUT(\mult_49/B_not [2]) );
  INV \mult_49/AN1_1_0  ( .IN(B[1]), .OUT(\mult_49/B_not [1]) );
  INV \mult_49/AN1_0_0  ( .IN(B[0]), .OUT(\mult_49/B_not [0]) );
  NOR2 \mult_49/AN3_31_0  ( .A(\mult_49/A_not [31]), .B(\mult_49/B_notx[0] ), 
        .OUT(\mult_49/ab[31][0] ) );
  NOR2 \mult_49/AN1_30_1  ( .A(\mult_49/A_not [30]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[30][1] ) );
  NOR2 \mult_49/AN1_30_0_0  ( .A(\mult_49/A_not [30]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[30][0] ) );
  NOR2 \mult_49/AN1_29_2  ( .A(\mult_49/A_not [29]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[29][2] ) );
  NOR2 \mult_49/AN1_29_1  ( .A(\mult_49/A_not [29]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[29][1] ) );
  NOR2 \mult_49/AN1_29_0_0  ( .A(\mult_49/A_not [29]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[29][0] ) );
  NOR2 \mult_49/AN1_28_3  ( .A(\mult_49/A_not [28]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[28][3] ) );
  NOR2 \mult_49/AN1_28_2  ( .A(\mult_49/A_not [28]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[28][2] ) );
  NOR2 \mult_49/AN1_28_1  ( .A(\mult_49/A_not [28]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[28][1] ) );
  NOR2 \mult_49/AN1_28_0_0  ( .A(\mult_49/A_not [28]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[28][0] ) );
  NOR2 \mult_49/AN1_27_4  ( .A(\mult_49/A_not [27]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[27][4] ) );
  NOR2 \mult_49/AN1_27_3  ( .A(\mult_49/A_not [27]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[27][3] ) );
  NOR2 \mult_49/AN1_27_2  ( .A(\mult_49/A_not [27]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[27][2] ) );
  NOR2 \mult_49/AN1_27_1  ( .A(\mult_49/A_not [27]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[27][1] ) );
  NOR2 \mult_49/AN1_27_0_0  ( .A(\mult_49/A_not [27]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[27][0] ) );
  NOR2 \mult_49/AN1_26_5  ( .A(\mult_49/A_not [26]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[26][5] ) );
  NOR2 \mult_49/AN1_26_4  ( .A(\mult_49/A_not [26]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[26][4] ) );
  NOR2 \mult_49/AN1_26_3  ( .A(\mult_49/A_not [26]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[26][3] ) );
  NOR2 \mult_49/AN1_26_2  ( .A(\mult_49/A_not [26]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[26][2] ) );
  NOR2 \mult_49/AN1_26_1  ( .A(\mult_49/A_not [26]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[26][1] ) );
  NOR2 \mult_49/AN1_26_0_0  ( .A(\mult_49/A_not [26]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[26][0] ) );
  NOR2 \mult_49/AN1_25_6  ( .A(\mult_49/A_not [25]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[25][6] ) );
  NOR2 \mult_49/AN1_25_5  ( .A(\mult_49/A_not [25]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[25][5] ) );
  NOR2 \mult_49/AN1_25_4  ( .A(\mult_49/A_not [25]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[25][4] ) );
  NOR2 \mult_49/AN1_25_3  ( .A(\mult_49/A_not [25]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[25][3] ) );
  NOR2 \mult_49/AN1_25_2  ( .A(\mult_49/A_not [25]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[25][2] ) );
  NOR2 \mult_49/AN1_25_1  ( .A(\mult_49/A_not [25]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[25][1] ) );
  NOR2 \mult_49/AN1_25_0_0  ( .A(\mult_49/A_not [25]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[25][0] ) );
  NOR2 \mult_49/AN1_24_7  ( .A(\mult_49/A_not [24]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[24][7] ) );
  NOR2 \mult_49/AN1_24_6  ( .A(\mult_49/A_not [24]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[24][6] ) );
  NOR2 \mult_49/AN1_24_5  ( .A(\mult_49/A_not [24]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[24][5] ) );
  NOR2 \mult_49/AN1_24_4  ( .A(\mult_49/A_not [24]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[24][4] ) );
  NOR2 \mult_49/AN1_24_3  ( .A(\mult_49/A_not [24]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[24][3] ) );
  NOR2 \mult_49/AN1_24_2  ( .A(\mult_49/A_not [24]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[24][2] ) );
  NOR2 \mult_49/AN1_24_1  ( .A(\mult_49/A_not [24]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[24][1] ) );
  NOR2 \mult_49/AN1_24_0_0  ( .A(\mult_49/A_not [24]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[24][0] ) );
  NOR2 \mult_49/AN1_23_8  ( .A(\mult_49/A_not [23]), .B(\mult_49/B_not [8]), 
        .OUT(\mult_49/ab[23][8] ) );
  NOR2 \mult_49/AN1_23_7  ( .A(\mult_49/A_not [23]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[23][7] ) );
  NOR2 \mult_49/AN1_23_6  ( .A(\mult_49/A_not [23]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[23][6] ) );
  NOR2 \mult_49/AN1_23_5  ( .A(\mult_49/A_not [23]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[23][5] ) );
  NOR2 \mult_49/AN1_23_4  ( .A(\mult_49/A_not [23]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[23][4] ) );
  NOR2 \mult_49/AN1_23_3  ( .A(\mult_49/A_not [23]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[23][3] ) );
  NOR2 \mult_49/AN1_23_2  ( .A(\mult_49/A_not [23]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[23][2] ) );
  NOR2 \mult_49/AN1_23_1  ( .A(\mult_49/A_not [23]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[23][1] ) );
  NOR2 \mult_49/AN1_23_0_0  ( .A(\mult_49/A_not [23]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[23][0] ) );
  NOR2 \mult_49/AN1_22_9  ( .A(\mult_49/A_not [22]), .B(\mult_49/B_not [9]), 
        .OUT(\mult_49/ab[22][9] ) );
  NOR2 \mult_49/AN1_22_8  ( .A(\mult_49/A_not [22]), .B(\mult_49/B_not [8]), 
        .OUT(\mult_49/ab[22][8] ) );
  NOR2 \mult_49/AN1_22_7  ( .A(\mult_49/A_not [22]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[22][7] ) );
  NOR2 \mult_49/AN1_22_6  ( .A(\mult_49/A_not [22]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[22][6] ) );
  NOR2 \mult_49/AN1_22_5  ( .A(\mult_49/A_not [22]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[22][5] ) );
  NOR2 \mult_49/AN1_22_4  ( .A(\mult_49/A_not [22]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[22][4] ) );
  NOR2 \mult_49/AN1_22_3  ( .A(\mult_49/A_not [22]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[22][3] ) );
  NOR2 \mult_49/AN1_22_2  ( .A(\mult_49/A_not [22]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[22][2] ) );
  NOR2 \mult_49/AN1_22_1  ( .A(\mult_49/A_not [22]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[22][1] ) );
  NOR2 \mult_49/AN1_22_0_0  ( .A(\mult_49/A_not [22]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[22][0] ) );
  NOR2 \mult_49/AN1_21_10  ( .A(\mult_49/A_not [21]), .B(\mult_49/B_not [10]), 
        .OUT(\mult_49/ab[21][10] ) );
  NOR2 \mult_49/AN1_21_9  ( .A(\mult_49/A_not [21]), .B(\mult_49/B_not [9]), 
        .OUT(\mult_49/ab[21][9] ) );
  NOR2 \mult_49/AN1_21_8  ( .A(\mult_49/A_not [21]), .B(\mult_49/B_not [8]), 
        .OUT(\mult_49/ab[21][8] ) );
  NOR2 \mult_49/AN1_21_7  ( .A(\mult_49/A_not [21]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[21][7] ) );
  NOR2 \mult_49/AN1_21_6  ( .A(\mult_49/A_not [21]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[21][6] ) );
  NOR2 \mult_49/AN1_21_5  ( .A(\mult_49/A_not [21]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[21][5] ) );
  NOR2 \mult_49/AN1_21_4  ( .A(\mult_49/A_not [21]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[21][4] ) );
  NOR2 \mult_49/AN1_21_3  ( .A(\mult_49/A_not [21]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[21][3] ) );
  NOR2 \mult_49/AN1_21_2  ( .A(\mult_49/A_not [21]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[21][2] ) );
  NOR2 \mult_49/AN1_21_1  ( .A(\mult_49/A_not [21]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[21][1] ) );
  NOR2 \mult_49/AN1_21_0_0  ( .A(\mult_49/A_not [21]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[21][0] ) );
  NOR2 \mult_49/AN1_20_11  ( .A(\mult_49/A_not [20]), .B(\mult_49/B_not [11]), 
        .OUT(\mult_49/ab[20][11] ) );
  NOR2 \mult_49/AN1_20_10  ( .A(\mult_49/A_not [20]), .B(\mult_49/B_not [10]), 
        .OUT(\mult_49/ab[20][10] ) );
  NOR2 \mult_49/AN1_20_9  ( .A(\mult_49/A_not [20]), .B(\mult_49/B_not [9]), 
        .OUT(\mult_49/ab[20][9] ) );
  NOR2 \mult_49/AN1_20_8  ( .A(\mult_49/A_not [20]), .B(\mult_49/B_not [8]), 
        .OUT(\mult_49/ab[20][8] ) );
  NOR2 \mult_49/AN1_20_7  ( .A(\mult_49/A_not [20]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[20][7] ) );
  NOR2 \mult_49/AN1_20_6  ( .A(\mult_49/A_not [20]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[20][6] ) );
  NOR2 \mult_49/AN1_20_5  ( .A(\mult_49/A_not [20]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[20][5] ) );
  NOR2 \mult_49/AN1_20_4  ( .A(\mult_49/A_not [20]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[20][4] ) );
  NOR2 \mult_49/AN1_20_3  ( .A(\mult_49/A_not [20]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[20][3] ) );
  NOR2 \mult_49/AN1_20_2  ( .A(\mult_49/A_not [20]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[20][2] ) );
  NOR2 \mult_49/AN1_20_1  ( .A(\mult_49/A_not [20]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[20][1] ) );
  NOR2 \mult_49/AN1_20_0_0  ( .A(\mult_49/A_not [20]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[20][0] ) );
  NOR2 \mult_49/AN1_19_12  ( .A(\mult_49/A_not [19]), .B(\mult_49/B_not [12]), 
        .OUT(\mult_49/ab[19][12] ) );
  NOR2 \mult_49/AN1_19_11  ( .A(\mult_49/A_not [19]), .B(\mult_49/B_not [11]), 
        .OUT(\mult_49/ab[19][11] ) );
  NOR2 \mult_49/AN1_19_10  ( .A(\mult_49/A_not [19]), .B(\mult_49/B_not [10]), 
        .OUT(\mult_49/ab[19][10] ) );
  NOR2 \mult_49/AN1_19_9  ( .A(\mult_49/A_not [19]), .B(\mult_49/B_not [9]), 
        .OUT(\mult_49/ab[19][9] ) );
  NOR2 \mult_49/AN1_19_8  ( .A(\mult_49/A_not [19]), .B(\mult_49/B_not [8]), 
        .OUT(\mult_49/ab[19][8] ) );
  NOR2 \mult_49/AN1_19_7  ( .A(\mult_49/A_not [19]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[19][7] ) );
  NOR2 \mult_49/AN1_19_6  ( .A(\mult_49/A_not [19]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[19][6] ) );
  NOR2 \mult_49/AN1_19_5  ( .A(\mult_49/A_not [19]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[19][5] ) );
  NOR2 \mult_49/AN1_19_4  ( .A(\mult_49/A_not [19]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[19][4] ) );
  NOR2 \mult_49/AN1_19_3  ( .A(\mult_49/A_not [19]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[19][3] ) );
  NOR2 \mult_49/AN1_19_2  ( .A(\mult_49/A_not [19]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[19][2] ) );
  NOR2 \mult_49/AN1_19_1  ( .A(\mult_49/A_not [19]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[19][1] ) );
  NOR2 \mult_49/AN1_19_0_0  ( .A(\mult_49/A_not [19]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[19][0] ) );
  NOR2 \mult_49/AN1_18_13  ( .A(\mult_49/A_not [18]), .B(\mult_49/B_not [13]), 
        .OUT(\mult_49/ab[18][13] ) );
  NOR2 \mult_49/AN1_18_12  ( .A(\mult_49/A_not [18]), .B(\mult_49/B_not [12]), 
        .OUT(\mult_49/ab[18][12] ) );
  NOR2 \mult_49/AN1_18_11  ( .A(\mult_49/A_not [18]), .B(\mult_49/B_not [11]), 
        .OUT(\mult_49/ab[18][11] ) );
  NOR2 \mult_49/AN1_18_10  ( .A(\mult_49/A_not [18]), .B(\mult_49/B_not [10]), 
        .OUT(\mult_49/ab[18][10] ) );
  NOR2 \mult_49/AN1_18_9  ( .A(\mult_49/A_not [18]), .B(\mult_49/B_not [9]), 
        .OUT(\mult_49/ab[18][9] ) );
  NOR2 \mult_49/AN1_18_8  ( .A(\mult_49/A_not [18]), .B(\mult_49/B_not [8]), 
        .OUT(\mult_49/ab[18][8] ) );
  NOR2 \mult_49/AN1_18_7  ( .A(\mult_49/A_not [18]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[18][7] ) );
  NOR2 \mult_49/AN1_18_6  ( .A(\mult_49/A_not [18]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[18][6] ) );
  NOR2 \mult_49/AN1_18_5  ( .A(\mult_49/A_not [18]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[18][5] ) );
  NOR2 \mult_49/AN1_18_4  ( .A(\mult_49/A_not [18]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[18][4] ) );
  NOR2 \mult_49/AN1_18_3  ( .A(\mult_49/A_not [18]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[18][3] ) );
  NOR2 \mult_49/AN1_18_2  ( .A(\mult_49/A_not [18]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[18][2] ) );
  NOR2 \mult_49/AN1_18_1  ( .A(\mult_49/A_not [18]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[18][1] ) );
  NOR2 \mult_49/AN1_18_0_0  ( .A(\mult_49/A_not [18]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[18][0] ) );
  NOR2 \mult_49/AN1_17_14  ( .A(\mult_49/A_not [17]), .B(\mult_49/B_not [14]), 
        .OUT(\mult_49/ab[17][14] ) );
  NOR2 \mult_49/AN1_17_13  ( .A(\mult_49/A_not [17]), .B(\mult_49/B_not [13]), 
        .OUT(\mult_49/ab[17][13] ) );
  NOR2 \mult_49/AN1_17_12  ( .A(\mult_49/A_not [17]), .B(\mult_49/B_not [12]), 
        .OUT(\mult_49/ab[17][12] ) );
  NOR2 \mult_49/AN1_17_11  ( .A(\mult_49/A_not [17]), .B(\mult_49/B_not [11]), 
        .OUT(\mult_49/ab[17][11] ) );
  NOR2 \mult_49/AN1_17_10  ( .A(\mult_49/A_not [17]), .B(\mult_49/B_not [10]), 
        .OUT(\mult_49/ab[17][10] ) );
  NOR2 \mult_49/AN1_17_9  ( .A(\mult_49/A_not [17]), .B(\mult_49/B_not [9]), 
        .OUT(\mult_49/ab[17][9] ) );
  NOR2 \mult_49/AN1_17_8  ( .A(\mult_49/A_not [17]), .B(\mult_49/B_not [8]), 
        .OUT(\mult_49/ab[17][8] ) );
  NOR2 \mult_49/AN1_17_7  ( .A(\mult_49/A_not [17]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[17][7] ) );
  NOR2 \mult_49/AN1_17_6  ( .A(\mult_49/A_not [17]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[17][6] ) );
  NOR2 \mult_49/AN1_17_5  ( .A(\mult_49/A_not [17]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[17][5] ) );
  NOR2 \mult_49/AN1_17_4  ( .A(\mult_49/A_not [17]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[17][4] ) );
  NOR2 \mult_49/AN1_17_3  ( .A(\mult_49/A_not [17]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[17][3] ) );
  NOR2 \mult_49/AN1_17_2  ( .A(\mult_49/A_not [17]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[17][2] ) );
  NOR2 \mult_49/AN1_17_1  ( .A(\mult_49/A_not [17]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[17][1] ) );
  NOR2 \mult_49/AN1_17_0_0  ( .A(\mult_49/A_not [17]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[17][0] ) );
  NOR2 \mult_49/AN1_16_15  ( .A(\mult_49/A_not [16]), .B(\mult_49/B_not [15]), 
        .OUT(\mult_49/ab[16][15] ) );
  NOR2 \mult_49/AN1_16_14  ( .A(\mult_49/A_not [16]), .B(\mult_49/B_not [14]), 
        .OUT(\mult_49/ab[16][14] ) );
  NOR2 \mult_49/AN1_16_13  ( .A(\mult_49/A_not [16]), .B(\mult_49/B_not [13]), 
        .OUT(\mult_49/ab[16][13] ) );
  NOR2 \mult_49/AN1_16_12  ( .A(\mult_49/A_not [16]), .B(\mult_49/B_not [12]), 
        .OUT(\mult_49/ab[16][12] ) );
  NOR2 \mult_49/AN1_16_11  ( .A(\mult_49/A_not [16]), .B(\mult_49/B_not [11]), 
        .OUT(\mult_49/ab[16][11] ) );
  NOR2 \mult_49/AN1_16_10  ( .A(\mult_49/A_not [16]), .B(\mult_49/B_not [10]), 
        .OUT(\mult_49/ab[16][10] ) );
  NOR2 \mult_49/AN1_16_9  ( .A(\mult_49/A_not [16]), .B(\mult_49/B_not [9]), 
        .OUT(\mult_49/ab[16][9] ) );
  NOR2 \mult_49/AN1_16_8  ( .A(\mult_49/A_not [16]), .B(\mult_49/B_not [8]), 
        .OUT(\mult_49/ab[16][8] ) );
  NOR2 \mult_49/AN1_16_7  ( .A(\mult_49/A_not [16]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[16][7] ) );
  NOR2 \mult_49/AN1_16_6  ( .A(\mult_49/A_not [16]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[16][6] ) );
  NOR2 \mult_49/AN1_16_5  ( .A(\mult_49/A_not [16]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[16][5] ) );
  NOR2 \mult_49/AN1_16_4  ( .A(\mult_49/A_not [16]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[16][4] ) );
  NOR2 \mult_49/AN1_16_3  ( .A(\mult_49/A_not [16]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[16][3] ) );
  NOR2 \mult_49/AN1_16_2  ( .A(\mult_49/A_not [16]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[16][2] ) );
  NOR2 \mult_49/AN1_16_1  ( .A(\mult_49/A_not [16]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[16][1] ) );
  NOR2 \mult_49/AN1_16_0_0  ( .A(\mult_49/A_not [16]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[16][0] ) );
  NOR2 \mult_49/AN1_15_16  ( .A(\mult_49/A_not [15]), .B(\mult_49/B_not [16]), 
        .OUT(\mult_49/ab[15][16] ) );
  NOR2 \mult_49/AN1_15_15  ( .A(\mult_49/A_not [15]), .B(\mult_49/B_not [15]), 
        .OUT(\mult_49/ab[15][15] ) );
  NOR2 \mult_49/AN1_15_14  ( .A(\mult_49/A_not [15]), .B(\mult_49/B_not [14]), 
        .OUT(\mult_49/ab[15][14] ) );
  NOR2 \mult_49/AN1_15_13  ( .A(\mult_49/A_not [15]), .B(\mult_49/B_not [13]), 
        .OUT(\mult_49/ab[15][13] ) );
  NOR2 \mult_49/AN1_15_12  ( .A(\mult_49/A_not [15]), .B(\mult_49/B_not [12]), 
        .OUT(\mult_49/ab[15][12] ) );
  NOR2 \mult_49/AN1_15_11  ( .A(\mult_49/A_not [15]), .B(\mult_49/B_not [11]), 
        .OUT(\mult_49/ab[15][11] ) );
  NOR2 \mult_49/AN1_15_10  ( .A(\mult_49/A_not [15]), .B(\mult_49/B_not [10]), 
        .OUT(\mult_49/ab[15][10] ) );
  NOR2 \mult_49/AN1_15_9  ( .A(\mult_49/A_not [15]), .B(\mult_49/B_not [9]), 
        .OUT(\mult_49/ab[15][9] ) );
  NOR2 \mult_49/AN1_15_8  ( .A(\mult_49/A_not [15]), .B(\mult_49/B_not [8]), 
        .OUT(\mult_49/ab[15][8] ) );
  NOR2 \mult_49/AN1_15_7  ( .A(\mult_49/A_not [15]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[15][7] ) );
  NOR2 \mult_49/AN1_15_6  ( .A(\mult_49/A_not [15]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[15][6] ) );
  NOR2 \mult_49/AN1_15_5  ( .A(\mult_49/A_not [15]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[15][5] ) );
  NOR2 \mult_49/AN1_15_4  ( .A(\mult_49/A_not [15]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[15][4] ) );
  NOR2 \mult_49/AN1_15_3  ( .A(\mult_49/A_not [15]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[15][3] ) );
  NOR2 \mult_49/AN1_15_2  ( .A(\mult_49/A_not [15]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[15][2] ) );
  NOR2 \mult_49/AN1_15_1  ( .A(\mult_49/A_not [15]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[15][1] ) );
  NOR2 \mult_49/AN1_15_0_0  ( .A(\mult_49/A_not [15]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[15][0] ) );
  NOR2 \mult_49/AN1_14_17  ( .A(\mult_49/A_not [14]), .B(\mult_49/B_not [17]), 
        .OUT(\mult_49/ab[14][17] ) );
  NOR2 \mult_49/AN1_14_16  ( .A(\mult_49/A_not [14]), .B(\mult_49/B_not [16]), 
        .OUT(\mult_49/ab[14][16] ) );
  NOR2 \mult_49/AN1_14_15  ( .A(\mult_49/A_not [14]), .B(\mult_49/B_not [15]), 
        .OUT(\mult_49/ab[14][15] ) );
  NOR2 \mult_49/AN1_14_14  ( .A(\mult_49/A_not [14]), .B(\mult_49/B_not [14]), 
        .OUT(\mult_49/ab[14][14] ) );
  NOR2 \mult_49/AN1_14_13  ( .A(\mult_49/A_not [14]), .B(\mult_49/B_not [13]), 
        .OUT(\mult_49/ab[14][13] ) );
  NOR2 \mult_49/AN1_14_12  ( .A(\mult_49/A_not [14]), .B(\mult_49/B_not [12]), 
        .OUT(\mult_49/ab[14][12] ) );
  NOR2 \mult_49/AN1_14_11  ( .A(\mult_49/A_not [14]), .B(\mult_49/B_not [11]), 
        .OUT(\mult_49/ab[14][11] ) );
  NOR2 \mult_49/AN1_14_10  ( .A(\mult_49/A_not [14]), .B(\mult_49/B_not [10]), 
        .OUT(\mult_49/ab[14][10] ) );
  NOR2 \mult_49/AN1_14_9  ( .A(\mult_49/A_not [14]), .B(\mult_49/B_not [9]), 
        .OUT(\mult_49/ab[14][9] ) );
  NOR2 \mult_49/AN1_14_8  ( .A(\mult_49/A_not [14]), .B(\mult_49/B_not [8]), 
        .OUT(\mult_49/ab[14][8] ) );
  NOR2 \mult_49/AN1_14_7  ( .A(\mult_49/A_not [14]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[14][7] ) );
  NOR2 \mult_49/AN1_14_6  ( .A(\mult_49/A_not [14]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[14][6] ) );
  NOR2 \mult_49/AN1_14_5  ( .A(\mult_49/A_not [14]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[14][5] ) );
  NOR2 \mult_49/AN1_14_4  ( .A(\mult_49/A_not [14]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[14][4] ) );
  NOR2 \mult_49/AN1_14_3  ( .A(\mult_49/A_not [14]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[14][3] ) );
  NOR2 \mult_49/AN1_14_2  ( .A(\mult_49/A_not [14]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[14][2] ) );
  NOR2 \mult_49/AN1_14_1  ( .A(\mult_49/A_not [14]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[14][1] ) );
  NOR2 \mult_49/AN1_14_0_0  ( .A(\mult_49/A_not [14]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[14][0] ) );
  NOR2 \mult_49/AN1_13_18  ( .A(\mult_49/A_not [13]), .B(\mult_49/B_not [18]), 
        .OUT(\mult_49/ab[13][18] ) );
  NOR2 \mult_49/AN1_13_17  ( .A(\mult_49/A_not [13]), .B(\mult_49/B_not [17]), 
        .OUT(\mult_49/ab[13][17] ) );
  NOR2 \mult_49/AN1_13_16  ( .A(\mult_49/A_not [13]), .B(\mult_49/B_not [16]), 
        .OUT(\mult_49/ab[13][16] ) );
  NOR2 \mult_49/AN1_13_15  ( .A(\mult_49/A_not [13]), .B(\mult_49/B_not [15]), 
        .OUT(\mult_49/ab[13][15] ) );
  NOR2 \mult_49/AN1_13_14  ( .A(\mult_49/A_not [13]), .B(\mult_49/B_not [14]), 
        .OUT(\mult_49/ab[13][14] ) );
  NOR2 \mult_49/AN1_13_13  ( .A(\mult_49/A_not [13]), .B(\mult_49/B_not [13]), 
        .OUT(\mult_49/ab[13][13] ) );
  NOR2 \mult_49/AN1_13_12  ( .A(\mult_49/A_not [13]), .B(\mult_49/B_not [12]), 
        .OUT(\mult_49/ab[13][12] ) );
  NOR2 \mult_49/AN1_13_11  ( .A(\mult_49/A_not [13]), .B(\mult_49/B_not [11]), 
        .OUT(\mult_49/ab[13][11] ) );
  NOR2 \mult_49/AN1_13_10  ( .A(\mult_49/A_not [13]), .B(\mult_49/B_not [10]), 
        .OUT(\mult_49/ab[13][10] ) );
  NOR2 \mult_49/AN1_13_9  ( .A(\mult_49/A_not [13]), .B(\mult_49/B_not [9]), 
        .OUT(\mult_49/ab[13][9] ) );
  NOR2 \mult_49/AN1_13_8  ( .A(\mult_49/A_not [13]), .B(\mult_49/B_not [8]), 
        .OUT(\mult_49/ab[13][8] ) );
  NOR2 \mult_49/AN1_13_7  ( .A(\mult_49/A_not [13]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[13][7] ) );
  NOR2 \mult_49/AN1_13_6  ( .A(\mult_49/A_not [13]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[13][6] ) );
  NOR2 \mult_49/AN1_13_5  ( .A(\mult_49/A_not [13]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[13][5] ) );
  NOR2 \mult_49/AN1_13_4  ( .A(\mult_49/A_not [13]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[13][4] ) );
  NOR2 \mult_49/AN1_13_3  ( .A(\mult_49/A_not [13]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[13][3] ) );
  NOR2 \mult_49/AN1_13_2  ( .A(\mult_49/A_not [13]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[13][2] ) );
  NOR2 \mult_49/AN1_13_1  ( .A(\mult_49/A_not [13]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[13][1] ) );
  NOR2 \mult_49/AN1_13_0_0  ( .A(\mult_49/A_not [13]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[13][0] ) );
  NOR2 \mult_49/AN1_12_19  ( .A(\mult_49/A_not [12]), .B(\mult_49/B_not [19]), 
        .OUT(\mult_49/ab[12][19] ) );
  NOR2 \mult_49/AN1_12_18  ( .A(\mult_49/A_not [12]), .B(\mult_49/B_not [18]), 
        .OUT(\mult_49/ab[12][18] ) );
  NOR2 \mult_49/AN1_12_17  ( .A(\mult_49/A_not [12]), .B(\mult_49/B_not [17]), 
        .OUT(\mult_49/ab[12][17] ) );
  NOR2 \mult_49/AN1_12_16  ( .A(\mult_49/A_not [12]), .B(\mult_49/B_not [16]), 
        .OUT(\mult_49/ab[12][16] ) );
  NOR2 \mult_49/AN1_12_15  ( .A(\mult_49/A_not [12]), .B(\mult_49/B_not [15]), 
        .OUT(\mult_49/ab[12][15] ) );
  NOR2 \mult_49/AN1_12_14  ( .A(\mult_49/A_not [12]), .B(\mult_49/B_not [14]), 
        .OUT(\mult_49/ab[12][14] ) );
  NOR2 \mult_49/AN1_12_13  ( .A(\mult_49/A_not [12]), .B(\mult_49/B_not [13]), 
        .OUT(\mult_49/ab[12][13] ) );
  NOR2 \mult_49/AN1_12_12  ( .A(\mult_49/A_not [12]), .B(\mult_49/B_not [12]), 
        .OUT(\mult_49/ab[12][12] ) );
  NOR2 \mult_49/AN1_12_11  ( .A(\mult_49/A_not [12]), .B(\mult_49/B_not [11]), 
        .OUT(\mult_49/ab[12][11] ) );
  NOR2 \mult_49/AN1_12_10  ( .A(\mult_49/A_not [12]), .B(\mult_49/B_not [10]), 
        .OUT(\mult_49/ab[12][10] ) );
  NOR2 \mult_49/AN1_12_9  ( .A(\mult_49/A_not [12]), .B(\mult_49/B_not [9]), 
        .OUT(\mult_49/ab[12][9] ) );
  NOR2 \mult_49/AN1_12_8  ( .A(\mult_49/A_not [12]), .B(\mult_49/B_not [8]), 
        .OUT(\mult_49/ab[12][8] ) );
  NOR2 \mult_49/AN1_12_7  ( .A(\mult_49/A_not [12]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[12][7] ) );
  NOR2 \mult_49/AN1_12_6  ( .A(\mult_49/A_not [12]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[12][6] ) );
  NOR2 \mult_49/AN1_12_5  ( .A(\mult_49/A_not [12]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[12][5] ) );
  NOR2 \mult_49/AN1_12_4  ( .A(\mult_49/A_not [12]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[12][4] ) );
  NOR2 \mult_49/AN1_12_3  ( .A(\mult_49/A_not [12]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[12][3] ) );
  NOR2 \mult_49/AN1_12_2  ( .A(\mult_49/A_not [12]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[12][2] ) );
  NOR2 \mult_49/AN1_12_1  ( .A(\mult_49/A_not [12]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[12][1] ) );
  NOR2 \mult_49/AN1_12_0_0  ( .A(\mult_49/A_not [12]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[12][0] ) );
  NOR2 \mult_49/AN1_11_20  ( .A(\mult_49/A_not [11]), .B(\mult_49/B_not [20]), 
        .OUT(\mult_49/ab[11][20] ) );
  NOR2 \mult_49/AN1_11_19  ( .A(\mult_49/A_not [11]), .B(\mult_49/B_not [19]), 
        .OUT(\mult_49/ab[11][19] ) );
  NOR2 \mult_49/AN1_11_18  ( .A(\mult_49/A_not [11]), .B(\mult_49/B_not [18]), 
        .OUT(\mult_49/ab[11][18] ) );
  NOR2 \mult_49/AN1_11_17  ( .A(\mult_49/A_not [11]), .B(\mult_49/B_not [17]), 
        .OUT(\mult_49/ab[11][17] ) );
  NOR2 \mult_49/AN1_11_16  ( .A(\mult_49/A_not [11]), .B(\mult_49/B_not [16]), 
        .OUT(\mult_49/ab[11][16] ) );
  NOR2 \mult_49/AN1_11_15  ( .A(\mult_49/A_not [11]), .B(\mult_49/B_not [15]), 
        .OUT(\mult_49/ab[11][15] ) );
  NOR2 \mult_49/AN1_11_14  ( .A(\mult_49/A_not [11]), .B(\mult_49/B_not [14]), 
        .OUT(\mult_49/ab[11][14] ) );
  NOR2 \mult_49/AN1_11_13  ( .A(\mult_49/A_not [11]), .B(\mult_49/B_not [13]), 
        .OUT(\mult_49/ab[11][13] ) );
  NOR2 \mult_49/AN1_11_12  ( .A(\mult_49/A_not [11]), .B(\mult_49/B_not [12]), 
        .OUT(\mult_49/ab[11][12] ) );
  NOR2 \mult_49/AN1_11_11  ( .A(\mult_49/A_not [11]), .B(\mult_49/B_not [11]), 
        .OUT(\mult_49/ab[11][11] ) );
  NOR2 \mult_49/AN1_11_10  ( .A(\mult_49/A_not [11]), .B(\mult_49/B_not [10]), 
        .OUT(\mult_49/ab[11][10] ) );
  NOR2 \mult_49/AN1_11_9  ( .A(\mult_49/A_not [11]), .B(\mult_49/B_not [9]), 
        .OUT(\mult_49/ab[11][9] ) );
  NOR2 \mult_49/AN1_11_8  ( .A(\mult_49/A_not [11]), .B(\mult_49/B_not [8]), 
        .OUT(\mult_49/ab[11][8] ) );
  NOR2 \mult_49/AN1_11_7  ( .A(\mult_49/A_not [11]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[11][7] ) );
  NOR2 \mult_49/AN1_11_6  ( .A(\mult_49/A_not [11]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[11][6] ) );
  NOR2 \mult_49/AN1_11_5  ( .A(\mult_49/A_not [11]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[11][5] ) );
  NOR2 \mult_49/AN1_11_4  ( .A(\mult_49/A_not [11]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[11][4] ) );
  NOR2 \mult_49/AN1_11_3  ( .A(\mult_49/A_not [11]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[11][3] ) );
  NOR2 \mult_49/AN1_11_2  ( .A(\mult_49/A_not [11]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[11][2] ) );
  NOR2 \mult_49/AN1_11_1  ( .A(\mult_49/A_not [11]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[11][1] ) );
  NOR2 \mult_49/AN1_11_0_0  ( .A(\mult_49/A_not [11]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[11][0] ) );
  NOR2 \mult_49/AN1_10_21  ( .A(\mult_49/A_not [10]), .B(\mult_49/B_not [21]), 
        .OUT(\mult_49/ab[10][21] ) );
  NOR2 \mult_49/AN1_10_20  ( .A(\mult_49/A_not [10]), .B(\mult_49/B_not [20]), 
        .OUT(\mult_49/ab[10][20] ) );
  NOR2 \mult_49/AN1_10_19  ( .A(\mult_49/A_not [10]), .B(\mult_49/B_not [19]), 
        .OUT(\mult_49/ab[10][19] ) );
  NOR2 \mult_49/AN1_10_18  ( .A(\mult_49/A_not [10]), .B(\mult_49/B_not [18]), 
        .OUT(\mult_49/ab[10][18] ) );
  NOR2 \mult_49/AN1_10_17  ( .A(\mult_49/A_not [10]), .B(\mult_49/B_not [17]), 
        .OUT(\mult_49/ab[10][17] ) );
  NOR2 \mult_49/AN1_10_16  ( .A(\mult_49/A_not [10]), .B(\mult_49/B_not [16]), 
        .OUT(\mult_49/ab[10][16] ) );
  NOR2 \mult_49/AN1_10_15  ( .A(\mult_49/A_not [10]), .B(\mult_49/B_not [15]), 
        .OUT(\mult_49/ab[10][15] ) );
  NOR2 \mult_49/AN1_10_14  ( .A(\mult_49/A_not [10]), .B(\mult_49/B_not [14]), 
        .OUT(\mult_49/ab[10][14] ) );
  NOR2 \mult_49/AN1_10_13  ( .A(\mult_49/A_not [10]), .B(\mult_49/B_not [13]), 
        .OUT(\mult_49/ab[10][13] ) );
  NOR2 \mult_49/AN1_10_12  ( .A(\mult_49/A_not [10]), .B(\mult_49/B_not [12]), 
        .OUT(\mult_49/ab[10][12] ) );
  NOR2 \mult_49/AN1_10_11  ( .A(\mult_49/A_not [10]), .B(\mult_49/B_not [11]), 
        .OUT(\mult_49/ab[10][11] ) );
  NOR2 \mult_49/AN1_10_10  ( .A(\mult_49/A_not [10]), .B(\mult_49/B_not [10]), 
        .OUT(\mult_49/ab[10][10] ) );
  NOR2 \mult_49/AN1_10_9  ( .A(\mult_49/A_not [10]), .B(\mult_49/B_not [9]), 
        .OUT(\mult_49/ab[10][9] ) );
  NOR2 \mult_49/AN1_10_8  ( .A(\mult_49/A_not [10]), .B(\mult_49/B_not [8]), 
        .OUT(\mult_49/ab[10][8] ) );
  NOR2 \mult_49/AN1_10_7  ( .A(\mult_49/A_not [10]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[10][7] ) );
  NOR2 \mult_49/AN1_10_6  ( .A(\mult_49/A_not [10]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[10][6] ) );
  NOR2 \mult_49/AN1_10_5  ( .A(\mult_49/A_not [10]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[10][5] ) );
  NOR2 \mult_49/AN1_10_4  ( .A(\mult_49/A_not [10]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[10][4] ) );
  NOR2 \mult_49/AN1_10_3  ( .A(\mult_49/A_not [10]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[10][3] ) );
  NOR2 \mult_49/AN1_10_2  ( .A(\mult_49/A_not [10]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[10][2] ) );
  NOR2 \mult_49/AN1_10_1  ( .A(\mult_49/A_not [10]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[10][1] ) );
  NOR2 \mult_49/AN1_10_0_0  ( .A(\mult_49/A_not [10]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[10][0] ) );
  NOR2 \mult_49/AN1_9_22  ( .A(\mult_49/A_not [9]), .B(\mult_49/B_not [22]), 
        .OUT(\mult_49/ab[9][22] ) );
  NOR2 \mult_49/AN1_9_21  ( .A(\mult_49/A_not [9]), .B(\mult_49/B_not [21]), 
        .OUT(\mult_49/ab[9][21] ) );
  NOR2 \mult_49/AN1_9_20  ( .A(\mult_49/A_not [9]), .B(\mult_49/B_not [20]), 
        .OUT(\mult_49/ab[9][20] ) );
  NOR2 \mult_49/AN1_9_19  ( .A(\mult_49/A_not [9]), .B(\mult_49/B_not [19]), 
        .OUT(\mult_49/ab[9][19] ) );
  NOR2 \mult_49/AN1_9_18  ( .A(\mult_49/A_not [9]), .B(\mult_49/B_not [18]), 
        .OUT(\mult_49/ab[9][18] ) );
  NOR2 \mult_49/AN1_9_17  ( .A(\mult_49/A_not [9]), .B(\mult_49/B_not [17]), 
        .OUT(\mult_49/ab[9][17] ) );
  NOR2 \mult_49/AN1_9_16  ( .A(\mult_49/A_not [9]), .B(\mult_49/B_not [16]), 
        .OUT(\mult_49/ab[9][16] ) );
  NOR2 \mult_49/AN1_9_15  ( .A(\mult_49/A_not [9]), .B(\mult_49/B_not [15]), 
        .OUT(\mult_49/ab[9][15] ) );
  NOR2 \mult_49/AN1_9_14  ( .A(\mult_49/A_not [9]), .B(\mult_49/B_not [14]), 
        .OUT(\mult_49/ab[9][14] ) );
  NOR2 \mult_49/AN1_9_13  ( .A(\mult_49/A_not [9]), .B(\mult_49/B_not [13]), 
        .OUT(\mult_49/ab[9][13] ) );
  NOR2 \mult_49/AN1_9_12  ( .A(\mult_49/A_not [9]), .B(\mult_49/B_not [12]), 
        .OUT(\mult_49/ab[9][12] ) );
  NOR2 \mult_49/AN1_9_11  ( .A(\mult_49/A_not [9]), .B(\mult_49/B_not [11]), 
        .OUT(\mult_49/ab[9][11] ) );
  NOR2 \mult_49/AN1_9_10  ( .A(\mult_49/A_not [9]), .B(\mult_49/B_not [10]), 
        .OUT(\mult_49/ab[9][10] ) );
  NOR2 \mult_49/AN1_9_9  ( .A(\mult_49/A_not [9]), .B(\mult_49/B_not [9]), 
        .OUT(\mult_49/ab[9][9] ) );
  NOR2 \mult_49/AN1_9_8  ( .A(\mult_49/A_not [9]), .B(\mult_49/B_not [8]), 
        .OUT(\mult_49/ab[9][8] ) );
  NOR2 \mult_49/AN1_9_7  ( .A(\mult_49/A_not [9]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[9][7] ) );
  NOR2 \mult_49/AN1_9_6  ( .A(\mult_49/A_not [9]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[9][6] ) );
  NOR2 \mult_49/AN1_9_5  ( .A(\mult_49/A_not [9]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[9][5] ) );
  NOR2 \mult_49/AN1_9_4  ( .A(\mult_49/A_not [9]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[9][4] ) );
  NOR2 \mult_49/AN1_9_3  ( .A(\mult_49/A_not [9]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[9][3] ) );
  NOR2 \mult_49/AN1_9_2  ( .A(\mult_49/A_not [9]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[9][2] ) );
  NOR2 \mult_49/AN1_9_1  ( .A(\mult_49/A_not [9]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[9][1] ) );
  NOR2 \mult_49/AN1_9_0_0  ( .A(\mult_49/A_not [9]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[9][0] ) );
  NOR2 \mult_49/AN1_8_23  ( .A(\mult_49/A_not [8]), .B(\mult_49/B_not [23]), 
        .OUT(\mult_49/ab[8][23] ) );
  NOR2 \mult_49/AN1_8_22  ( .A(\mult_49/A_not [8]), .B(\mult_49/B_not [22]), 
        .OUT(\mult_49/ab[8][22] ) );
  NOR2 \mult_49/AN1_8_21  ( .A(\mult_49/A_not [8]), .B(\mult_49/B_not [21]), 
        .OUT(\mult_49/ab[8][21] ) );
  NOR2 \mult_49/AN1_8_20  ( .A(\mult_49/A_not [8]), .B(\mult_49/B_not [20]), 
        .OUT(\mult_49/ab[8][20] ) );
  NOR2 \mult_49/AN1_8_19  ( .A(\mult_49/A_not [8]), .B(\mult_49/B_not [19]), 
        .OUT(\mult_49/ab[8][19] ) );
  NOR2 \mult_49/AN1_8_18  ( .A(\mult_49/A_not [8]), .B(\mult_49/B_not [18]), 
        .OUT(\mult_49/ab[8][18] ) );
  NOR2 \mult_49/AN1_8_17  ( .A(\mult_49/A_not [8]), .B(\mult_49/B_not [17]), 
        .OUT(\mult_49/ab[8][17] ) );
  NOR2 \mult_49/AN1_8_16  ( .A(\mult_49/A_not [8]), .B(\mult_49/B_not [16]), 
        .OUT(\mult_49/ab[8][16] ) );
  NOR2 \mult_49/AN1_8_15  ( .A(\mult_49/A_not [8]), .B(\mult_49/B_not [15]), 
        .OUT(\mult_49/ab[8][15] ) );
  NOR2 \mult_49/AN1_8_14  ( .A(\mult_49/A_not [8]), .B(\mult_49/B_not [14]), 
        .OUT(\mult_49/ab[8][14] ) );
  NOR2 \mult_49/AN1_8_13  ( .A(\mult_49/A_not [8]), .B(\mult_49/B_not [13]), 
        .OUT(\mult_49/ab[8][13] ) );
  NOR2 \mult_49/AN1_8_12  ( .A(\mult_49/A_not [8]), .B(\mult_49/B_not [12]), 
        .OUT(\mult_49/ab[8][12] ) );
  NOR2 \mult_49/AN1_8_11  ( .A(\mult_49/A_not [8]), .B(\mult_49/B_not [11]), 
        .OUT(\mult_49/ab[8][11] ) );
  NOR2 \mult_49/AN1_8_10  ( .A(\mult_49/A_not [8]), .B(\mult_49/B_not [10]), 
        .OUT(\mult_49/ab[8][10] ) );
  NOR2 \mult_49/AN1_8_9  ( .A(\mult_49/A_not [8]), .B(\mult_49/B_not [9]), 
        .OUT(\mult_49/ab[8][9] ) );
  NOR2 \mult_49/AN1_8_8  ( .A(\mult_49/A_not [8]), .B(\mult_49/B_not [8]), 
        .OUT(\mult_49/ab[8][8] ) );
  NOR2 \mult_49/AN1_8_7  ( .A(\mult_49/A_not [8]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[8][7] ) );
  NOR2 \mult_49/AN1_8_6  ( .A(\mult_49/A_not [8]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[8][6] ) );
  NOR2 \mult_49/AN1_8_5  ( .A(\mult_49/A_not [8]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[8][5] ) );
  NOR2 \mult_49/AN1_8_4  ( .A(\mult_49/A_not [8]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[8][4] ) );
  NOR2 \mult_49/AN1_8_3  ( .A(\mult_49/A_not [8]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[8][3] ) );
  NOR2 \mult_49/AN1_8_2  ( .A(\mult_49/A_not [8]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[8][2] ) );
  NOR2 \mult_49/AN1_8_1  ( .A(\mult_49/A_not [8]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[8][1] ) );
  NOR2 \mult_49/AN1_8_0_0  ( .A(\mult_49/A_not [8]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[8][0] ) );
  NOR2 \mult_49/AN1_7_24  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [24]), 
        .OUT(\mult_49/ab[7][24] ) );
  NOR2 \mult_49/AN1_7_23  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [23]), 
        .OUT(\mult_49/ab[7][23] ) );
  NOR2 \mult_49/AN1_7_22  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [22]), 
        .OUT(\mult_49/ab[7][22] ) );
  NOR2 \mult_49/AN1_7_21  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [21]), 
        .OUT(\mult_49/ab[7][21] ) );
  NOR2 \mult_49/AN1_7_20  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [20]), 
        .OUT(\mult_49/ab[7][20] ) );
  NOR2 \mult_49/AN1_7_19  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [19]), 
        .OUT(\mult_49/ab[7][19] ) );
  NOR2 \mult_49/AN1_7_18  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [18]), 
        .OUT(\mult_49/ab[7][18] ) );
  NOR2 \mult_49/AN1_7_17  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [17]), 
        .OUT(\mult_49/ab[7][17] ) );
  NOR2 \mult_49/AN1_7_16  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [16]), 
        .OUT(\mult_49/ab[7][16] ) );
  NOR2 \mult_49/AN1_7_15  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [15]), 
        .OUT(\mult_49/ab[7][15] ) );
  NOR2 \mult_49/AN1_7_14  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [14]), 
        .OUT(\mult_49/ab[7][14] ) );
  NOR2 \mult_49/AN1_7_13  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [13]), 
        .OUT(\mult_49/ab[7][13] ) );
  NOR2 \mult_49/AN1_7_12  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [12]), 
        .OUT(\mult_49/ab[7][12] ) );
  NOR2 \mult_49/AN1_7_11  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [11]), 
        .OUT(\mult_49/ab[7][11] ) );
  NOR2 \mult_49/AN1_7_10  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [10]), 
        .OUT(\mult_49/ab[7][10] ) );
  NOR2 \mult_49/AN1_7_9  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [9]), 
        .OUT(\mult_49/ab[7][9] ) );
  NOR2 \mult_49/AN1_7_8  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [8]), 
        .OUT(\mult_49/ab[7][8] ) );
  NOR2 \mult_49/AN1_7_7  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[7][7] ) );
  NOR2 \mult_49/AN1_7_6  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[7][6] ) );
  NOR2 \mult_49/AN1_7_5  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[7][5] ) );
  NOR2 \mult_49/AN1_7_4  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[7][4] ) );
  NOR2 \mult_49/AN1_7_3  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[7][3] ) );
  NOR2 \mult_49/AN1_7_2  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[7][2] ) );
  NOR2 \mult_49/AN1_7_1  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[7][1] ) );
  NOR2 \mult_49/AN1_7_0_0  ( .A(\mult_49/A_not [7]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[7][0] ) );
  NOR2 \mult_49/AN1_6_25  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [25]), 
        .OUT(\mult_49/ab[6][25] ) );
  NOR2 \mult_49/AN1_6_24  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [24]), 
        .OUT(\mult_49/ab[6][24] ) );
  NOR2 \mult_49/AN1_6_23  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [23]), 
        .OUT(\mult_49/ab[6][23] ) );
  NOR2 \mult_49/AN1_6_22  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [22]), 
        .OUT(\mult_49/ab[6][22] ) );
  NOR2 \mult_49/AN1_6_21  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [21]), 
        .OUT(\mult_49/ab[6][21] ) );
  NOR2 \mult_49/AN1_6_20  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [20]), 
        .OUT(\mult_49/ab[6][20] ) );
  NOR2 \mult_49/AN1_6_19  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [19]), 
        .OUT(\mult_49/ab[6][19] ) );
  NOR2 \mult_49/AN1_6_18  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [18]), 
        .OUT(\mult_49/ab[6][18] ) );
  NOR2 \mult_49/AN1_6_17  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [17]), 
        .OUT(\mult_49/ab[6][17] ) );
  NOR2 \mult_49/AN1_6_16  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [16]), 
        .OUT(\mult_49/ab[6][16] ) );
  NOR2 \mult_49/AN1_6_15  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [15]), 
        .OUT(\mult_49/ab[6][15] ) );
  NOR2 \mult_49/AN1_6_14  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [14]), 
        .OUT(\mult_49/ab[6][14] ) );
  NOR2 \mult_49/AN1_6_13  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [13]), 
        .OUT(\mult_49/ab[6][13] ) );
  NOR2 \mult_49/AN1_6_12  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [12]), 
        .OUT(\mult_49/ab[6][12] ) );
  NOR2 \mult_49/AN1_6_11  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [11]), 
        .OUT(\mult_49/ab[6][11] ) );
  NOR2 \mult_49/AN1_6_10  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [10]), 
        .OUT(\mult_49/ab[6][10] ) );
  NOR2 \mult_49/AN1_6_9  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [9]), 
        .OUT(\mult_49/ab[6][9] ) );
  NOR2 \mult_49/AN1_6_8  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [8]), 
        .OUT(\mult_49/ab[6][8] ) );
  NOR2 \mult_49/AN1_6_7  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[6][7] ) );
  NOR2 \mult_49/AN1_6_6  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[6][6] ) );
  NOR2 \mult_49/AN1_6_5  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[6][5] ) );
  NOR2 \mult_49/AN1_6_4  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[6][4] ) );
  NOR2 \mult_49/AN1_6_3  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[6][3] ) );
  NOR2 \mult_49/AN1_6_2  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[6][2] ) );
  NOR2 \mult_49/AN1_6_1  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[6][1] ) );
  NOR2 \mult_49/AN1_6_0_0  ( .A(\mult_49/A_not [6]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[6][0] ) );
  NOR2 \mult_49/AN1_5_26  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [26]), 
        .OUT(\mult_49/ab[5][26] ) );
  NOR2 \mult_49/AN1_5_25  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [25]), 
        .OUT(\mult_49/ab[5][25] ) );
  NOR2 \mult_49/AN1_5_24  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [24]), 
        .OUT(\mult_49/ab[5][24] ) );
  NOR2 \mult_49/AN1_5_23  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [23]), 
        .OUT(\mult_49/ab[5][23] ) );
  NOR2 \mult_49/AN1_5_22  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [22]), 
        .OUT(\mult_49/ab[5][22] ) );
  NOR2 \mult_49/AN1_5_21  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [21]), 
        .OUT(\mult_49/ab[5][21] ) );
  NOR2 \mult_49/AN1_5_20  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [20]), 
        .OUT(\mult_49/ab[5][20] ) );
  NOR2 \mult_49/AN1_5_19  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [19]), 
        .OUT(\mult_49/ab[5][19] ) );
  NOR2 \mult_49/AN1_5_18  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [18]), 
        .OUT(\mult_49/ab[5][18] ) );
  NOR2 \mult_49/AN1_5_17  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [17]), 
        .OUT(\mult_49/ab[5][17] ) );
  NOR2 \mult_49/AN1_5_16  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [16]), 
        .OUT(\mult_49/ab[5][16] ) );
  NOR2 \mult_49/AN1_5_15  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [15]), 
        .OUT(\mult_49/ab[5][15] ) );
  NOR2 \mult_49/AN1_5_14  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [14]), 
        .OUT(\mult_49/ab[5][14] ) );
  NOR2 \mult_49/AN1_5_13  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [13]), 
        .OUT(\mult_49/ab[5][13] ) );
  NOR2 \mult_49/AN1_5_12  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [12]), 
        .OUT(\mult_49/ab[5][12] ) );
  NOR2 \mult_49/AN1_5_11  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [11]), 
        .OUT(\mult_49/ab[5][11] ) );
  NOR2 \mult_49/AN1_5_10  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [10]), 
        .OUT(\mult_49/ab[5][10] ) );
  NOR2 \mult_49/AN1_5_9  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [9]), 
        .OUT(\mult_49/ab[5][9] ) );
  NOR2 \mult_49/AN1_5_8  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [8]), 
        .OUT(\mult_49/ab[5][8] ) );
  NOR2 \mult_49/AN1_5_7  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[5][7] ) );
  NOR2 \mult_49/AN1_5_6  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[5][6] ) );
  NOR2 \mult_49/AN1_5_5  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[5][5] ) );
  NOR2 \mult_49/AN1_5_4  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[5][4] ) );
  NOR2 \mult_49/AN1_5_3  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[5][3] ) );
  NOR2 \mult_49/AN1_5_2  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[5][2] ) );
  NOR2 \mult_49/AN1_5_1  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[5][1] ) );
  NOR2 \mult_49/AN1_5_0_0  ( .A(\mult_49/A_not [5]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[5][0] ) );
  NOR2 \mult_49/AN1_4_27  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [27]), 
        .OUT(\mult_49/ab[4][27] ) );
  NOR2 \mult_49/AN1_4_26  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [26]), 
        .OUT(\mult_49/ab[4][26] ) );
  NOR2 \mult_49/AN1_4_25  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [25]), 
        .OUT(\mult_49/ab[4][25] ) );
  NOR2 \mult_49/AN1_4_24  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [24]), 
        .OUT(\mult_49/ab[4][24] ) );
  NOR2 \mult_49/AN1_4_23  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [23]), 
        .OUT(\mult_49/ab[4][23] ) );
  NOR2 \mult_49/AN1_4_22  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [22]), 
        .OUT(\mult_49/ab[4][22] ) );
  NOR2 \mult_49/AN1_4_21  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [21]), 
        .OUT(\mult_49/ab[4][21] ) );
  NOR2 \mult_49/AN1_4_20  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [20]), 
        .OUT(\mult_49/ab[4][20] ) );
  NOR2 \mult_49/AN1_4_19  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [19]), 
        .OUT(\mult_49/ab[4][19] ) );
  NOR2 \mult_49/AN1_4_18  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [18]), 
        .OUT(\mult_49/ab[4][18] ) );
  NOR2 \mult_49/AN1_4_17  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [17]), 
        .OUT(\mult_49/ab[4][17] ) );
  NOR2 \mult_49/AN1_4_16  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [16]), 
        .OUT(\mult_49/ab[4][16] ) );
  NOR2 \mult_49/AN1_4_15  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [15]), 
        .OUT(\mult_49/ab[4][15] ) );
  NOR2 \mult_49/AN1_4_14  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [14]), 
        .OUT(\mult_49/ab[4][14] ) );
  NOR2 \mult_49/AN1_4_13  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [13]), 
        .OUT(\mult_49/ab[4][13] ) );
  NOR2 \mult_49/AN1_4_12  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [12]), 
        .OUT(\mult_49/ab[4][12] ) );
  NOR2 \mult_49/AN1_4_11  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [11]), 
        .OUT(\mult_49/ab[4][11] ) );
  NOR2 \mult_49/AN1_4_10  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [10]), 
        .OUT(\mult_49/ab[4][10] ) );
  NOR2 \mult_49/AN1_4_9  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [9]), 
        .OUT(\mult_49/ab[4][9] ) );
  NOR2 \mult_49/AN1_4_8  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [8]), 
        .OUT(\mult_49/ab[4][8] ) );
  NOR2 \mult_49/AN1_4_7  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[4][7] ) );
  NOR2 \mult_49/AN1_4_6  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[4][6] ) );
  NOR2 \mult_49/AN1_4_5  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[4][5] ) );
  NOR2 \mult_49/AN1_4_4  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[4][4] ) );
  NOR2 \mult_49/AN1_4_3  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[4][3] ) );
  NOR2 \mult_49/AN1_4_2  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[4][2] ) );
  NOR2 \mult_49/AN1_4_1  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[4][1] ) );
  NOR2 \mult_49/AN1_4_0_0  ( .A(\mult_49/A_not [4]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[4][0] ) );
  NOR2 \mult_49/AN1_3_28  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [28]), 
        .OUT(\mult_49/ab[3][28] ) );
  NOR2 \mult_49/AN1_3_27  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [27]), 
        .OUT(\mult_49/ab[3][27] ) );
  NOR2 \mult_49/AN1_3_26  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [26]), 
        .OUT(\mult_49/ab[3][26] ) );
  NOR2 \mult_49/AN1_3_25  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [25]), 
        .OUT(\mult_49/ab[3][25] ) );
  NOR2 \mult_49/AN1_3_24  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [24]), 
        .OUT(\mult_49/ab[3][24] ) );
  NOR2 \mult_49/AN1_3_23  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [23]), 
        .OUT(\mult_49/ab[3][23] ) );
  NOR2 \mult_49/AN1_3_22  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [22]), 
        .OUT(\mult_49/ab[3][22] ) );
  NOR2 \mult_49/AN1_3_21  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [21]), 
        .OUT(\mult_49/ab[3][21] ) );
  NOR2 \mult_49/AN1_3_20  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [20]), 
        .OUT(\mult_49/ab[3][20] ) );
  NOR2 \mult_49/AN1_3_19  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [19]), 
        .OUT(\mult_49/ab[3][19] ) );
  NOR2 \mult_49/AN1_3_18  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [18]), 
        .OUT(\mult_49/ab[3][18] ) );
  NOR2 \mult_49/AN1_3_17  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [17]), 
        .OUT(\mult_49/ab[3][17] ) );
  NOR2 \mult_49/AN1_3_16  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [16]), 
        .OUT(\mult_49/ab[3][16] ) );
  NOR2 \mult_49/AN1_3_15  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [15]), 
        .OUT(\mult_49/ab[3][15] ) );
  NOR2 \mult_49/AN1_3_14  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [14]), 
        .OUT(\mult_49/ab[3][14] ) );
  NOR2 \mult_49/AN1_3_13  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [13]), 
        .OUT(\mult_49/ab[3][13] ) );
  NOR2 \mult_49/AN1_3_12  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [12]), 
        .OUT(\mult_49/ab[3][12] ) );
  NOR2 \mult_49/AN1_3_11  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [11]), 
        .OUT(\mult_49/ab[3][11] ) );
  NOR2 \mult_49/AN1_3_10  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [10]), 
        .OUT(\mult_49/ab[3][10] ) );
  NOR2 \mult_49/AN1_3_9  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [9]), 
        .OUT(\mult_49/ab[3][9] ) );
  NOR2 \mult_49/AN1_3_8  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [8]), 
        .OUT(\mult_49/ab[3][8] ) );
  NOR2 \mult_49/AN1_3_7  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[3][7] ) );
  NOR2 \mult_49/AN1_3_6  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[3][6] ) );
  NOR2 \mult_49/AN1_3_5  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[3][5] ) );
  NOR2 \mult_49/AN1_3_4  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[3][4] ) );
  NOR2 \mult_49/AN1_3_3  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[3][3] ) );
  NOR2 \mult_49/AN1_3_2  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[3][2] ) );
  NOR2 \mult_49/AN1_3_1  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[3][1] ) );
  NOR2 \mult_49/AN1_3_0_0  ( .A(\mult_49/A_not [3]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[3][0] ) );
  NOR2 \mult_49/AN1_2_29  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [29]), 
        .OUT(\mult_49/ab[2][29] ) );
  NOR2 \mult_49/AN1_2_28  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [28]), 
        .OUT(\mult_49/ab[2][28] ) );
  NOR2 \mult_49/AN1_2_27  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [27]), 
        .OUT(\mult_49/ab[2][27] ) );
  NOR2 \mult_49/AN1_2_26  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [26]), 
        .OUT(\mult_49/ab[2][26] ) );
  NOR2 \mult_49/AN1_2_25  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [25]), 
        .OUT(\mult_49/ab[2][25] ) );
  NOR2 \mult_49/AN1_2_24  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [24]), 
        .OUT(\mult_49/ab[2][24] ) );
  NOR2 \mult_49/AN1_2_23  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [23]), 
        .OUT(\mult_49/ab[2][23] ) );
  NOR2 \mult_49/AN1_2_22  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [22]), 
        .OUT(\mult_49/ab[2][22] ) );
  NOR2 \mult_49/AN1_2_21  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [21]), 
        .OUT(\mult_49/ab[2][21] ) );
  NOR2 \mult_49/AN1_2_20  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [20]), 
        .OUT(\mult_49/ab[2][20] ) );
  NOR2 \mult_49/AN1_2_19  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [19]), 
        .OUT(\mult_49/ab[2][19] ) );
  NOR2 \mult_49/AN1_2_18  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [18]), 
        .OUT(\mult_49/ab[2][18] ) );
  NOR2 \mult_49/AN1_2_17  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [17]), 
        .OUT(\mult_49/ab[2][17] ) );
  NOR2 \mult_49/AN1_2_16  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [16]), 
        .OUT(\mult_49/ab[2][16] ) );
  NOR2 \mult_49/AN1_2_15  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [15]), 
        .OUT(\mult_49/ab[2][15] ) );
  NOR2 \mult_49/AN1_2_14  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [14]), 
        .OUT(\mult_49/ab[2][14] ) );
  NOR2 \mult_49/AN1_2_13  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [13]), 
        .OUT(\mult_49/ab[2][13] ) );
  NOR2 \mult_49/AN1_2_12  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [12]), 
        .OUT(\mult_49/ab[2][12] ) );
  NOR2 \mult_49/AN1_2_11  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [11]), 
        .OUT(\mult_49/ab[2][11] ) );
  NOR2 \mult_49/AN1_2_10  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [10]), 
        .OUT(\mult_49/ab[2][10] ) );
  NOR2 \mult_49/AN1_2_9  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [9]), 
        .OUT(\mult_49/ab[2][9] ) );
  NOR2 \mult_49/AN1_2_8  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [8]), 
        .OUT(\mult_49/ab[2][8] ) );
  NOR2 \mult_49/AN1_2_7  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[2][7] ) );
  NOR2 \mult_49/AN1_2_6  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[2][6] ) );
  NOR2 \mult_49/AN1_2_5  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[2][5] ) );
  NOR2 \mult_49/AN1_2_4  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[2][4] ) );
  NOR2 \mult_49/AN1_2_3  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[2][3] ) );
  NOR2 \mult_49/AN1_2_2  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[2][2] ) );
  NOR2 \mult_49/AN1_2_1  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[2][1] ) );
  NOR2 \mult_49/AN1_2_0_0  ( .A(\mult_49/A_not [2]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[2][0] ) );
  NOR2 \mult_49/AN1_1_30  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [30]), 
        .OUT(\mult_49/ab[1][30] ) );
  NOR2 \mult_49/AN1_1_29  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [29]), 
        .OUT(\mult_49/ab[1][29] ) );
  NOR2 \mult_49/AN1_1_28  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [28]), 
        .OUT(\mult_49/ab[1][28] ) );
  NOR2 \mult_49/AN1_1_27  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [27]), 
        .OUT(\mult_49/ab[1][27] ) );
  NOR2 \mult_49/AN1_1_26  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [26]), 
        .OUT(\mult_49/ab[1][26] ) );
  NOR2 \mult_49/AN1_1_25  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [25]), 
        .OUT(\mult_49/ab[1][25] ) );
  NOR2 \mult_49/AN1_1_24  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [24]), 
        .OUT(\mult_49/ab[1][24] ) );
  NOR2 \mult_49/AN1_1_23  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [23]), 
        .OUT(\mult_49/ab[1][23] ) );
  NOR2 \mult_49/AN1_1_22  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [22]), 
        .OUT(\mult_49/ab[1][22] ) );
  NOR2 \mult_49/AN1_1_21  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [21]), 
        .OUT(\mult_49/ab[1][21] ) );
  NOR2 \mult_49/AN1_1_20  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [20]), 
        .OUT(\mult_49/ab[1][20] ) );
  NOR2 \mult_49/AN1_1_19  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [19]), 
        .OUT(\mult_49/ab[1][19] ) );
  NOR2 \mult_49/AN1_1_18  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [18]), 
        .OUT(\mult_49/ab[1][18] ) );
  NOR2 \mult_49/AN1_1_17  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [17]), 
        .OUT(\mult_49/ab[1][17] ) );
  NOR2 \mult_49/AN1_1_16  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [16]), 
        .OUT(\mult_49/ab[1][16] ) );
  NOR2 \mult_49/AN1_1_15  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [15]), 
        .OUT(\mult_49/ab[1][15] ) );
  NOR2 \mult_49/AN1_1_14  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [14]), 
        .OUT(\mult_49/ab[1][14] ) );
  NOR2 \mult_49/AN1_1_13  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [13]), 
        .OUT(\mult_49/ab[1][13] ) );
  NOR2 \mult_49/AN1_1_12  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [12]), 
        .OUT(\mult_49/ab[1][12] ) );
  NOR2 \mult_49/AN1_1_11  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [11]), 
        .OUT(\mult_49/ab[1][11] ) );
  NOR2 \mult_49/AN1_1_10  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [10]), 
        .OUT(\mult_49/ab[1][10] ) );
  NOR2 \mult_49/AN1_1_9  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [9]), 
        .OUT(\mult_49/ab[1][9] ) );
  NOR2 \mult_49/AN1_1_8  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [8]), 
        .OUT(\mult_49/ab[1][8] ) );
  NOR2 \mult_49/AN1_1_7  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[1][7] ) );
  NOR2 \mult_49/AN1_1_6  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[1][6] ) );
  NOR2 \mult_49/AN1_1_5  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[1][5] ) );
  NOR2 \mult_49/AN1_1_4  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[1][4] ) );
  NOR2 \mult_49/AN1_1_3  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[1][3] ) );
  NOR2 \mult_49/AN1_1_2  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[1][2] ) );
  NOR2 \mult_49/AN1_1_1  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[1][1] ) );
  NOR2 \mult_49/AN1_1_0_0  ( .A(\mult_49/A_not [1]), .B(\mult_49/B_not [0]), 
        .OUT(\mult_49/ab[1][0] ) );
  NOR2 \mult_49/AN2_0_31  ( .A(\mult_49/A_notx[0] ), .B(\mult_49/B_not [31]), 
        .OUT(\mult_49/ab[0][31] ) );
  NOR2 \mult_49/AN1_0_30  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [30]), 
        .OUT(\mult_49/ab[0][30] ) );
  NOR2 \mult_49/AN1_0_29  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [29]), 
        .OUT(\mult_49/ab[0][29] ) );
  NOR2 \mult_49/AN1_0_28  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [28]), 
        .OUT(\mult_49/ab[0][28] ) );
  NOR2 \mult_49/AN1_0_27  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [27]), 
        .OUT(\mult_49/ab[0][27] ) );
  NOR2 \mult_49/AN1_0_26  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [26]), 
        .OUT(\mult_49/ab[0][26] ) );
  NOR2 \mult_49/AN1_0_25  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [25]), 
        .OUT(\mult_49/ab[0][25] ) );
  NOR2 \mult_49/AN1_0_24  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [24]), 
        .OUT(\mult_49/ab[0][24] ) );
  NOR2 \mult_49/AN1_0_23  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [23]), 
        .OUT(\mult_49/ab[0][23] ) );
  NOR2 \mult_49/AN1_0_22  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [22]), 
        .OUT(\mult_49/ab[0][22] ) );
  NOR2 \mult_49/AN1_0_21  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [21]), 
        .OUT(\mult_49/ab[0][21] ) );
  NOR2 \mult_49/AN1_0_20  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [20]), 
        .OUT(\mult_49/ab[0][20] ) );
  NOR2 \mult_49/AN1_0_19  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [19]), 
        .OUT(\mult_49/ab[0][19] ) );
  NOR2 \mult_49/AN1_0_18  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [18]), 
        .OUT(\mult_49/ab[0][18] ) );
  NOR2 \mult_49/AN1_0_17  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [17]), 
        .OUT(\mult_49/ab[0][17] ) );
  NOR2 \mult_49/AN1_0_16  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [16]), 
        .OUT(\mult_49/ab[0][16] ) );
  NOR2 \mult_49/AN1_0_15  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [15]), 
        .OUT(\mult_49/ab[0][15] ) );
  NOR2 \mult_49/AN1_0_14  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [14]), 
        .OUT(\mult_49/ab[0][14] ) );
  NOR2 \mult_49/AN1_0_13  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [13]), 
        .OUT(\mult_49/ab[0][13] ) );
  NOR2 \mult_49/AN1_0_12  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [12]), 
        .OUT(\mult_49/ab[0][12] ) );
  NOR2 \mult_49/AN1_0_11  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [11]), 
        .OUT(\mult_49/ab[0][11] ) );
  NOR2 \mult_49/AN1_0_10  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [10]), 
        .OUT(\mult_49/ab[0][10] ) );
  NOR2 \mult_49/AN1_0_9  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [9]), 
        .OUT(\mult_49/ab[0][9] ) );
  NOR2 \mult_49/AN1_0_8  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [8]), 
        .OUT(\mult_49/ab[0][8] ) );
  NOR2 \mult_49/AN1_0_7  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [7]), 
        .OUT(\mult_49/ab[0][7] ) );
  NOR2 \mult_49/AN1_0_6  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [6]), 
        .OUT(\mult_49/ab[0][6] ) );
  NOR2 \mult_49/AN1_0_5  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [5]), 
        .OUT(\mult_49/ab[0][5] ) );
  NOR2 \mult_49/AN1_0_4  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [4]), 
        .OUT(\mult_49/ab[0][4] ) );
  NOR2 \mult_49/AN1_0_3  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [3]), 
        .OUT(\mult_49/ab[0][3] ) );
  NOR2 \mult_49/AN1_0_2  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [2]), 
        .OUT(\mult_49/ab[0][2] ) );
  NOR2 \mult_49/AN1_0_1  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [1]), 
        .OUT(\mult_49/ab[0][1] ) );
  NOR2 \mult_49/AN1_0_0_0  ( .A(\mult_49/A_not [0]), .B(\mult_49/B_not [0]), 
        .OUT(N222) );
  NOR2 \gt_48/ULTI0_0  ( .A(B[0]), .B(n6462), .OUT(n6461) );
  NOR2 \gt_48/ULTI0_1  ( .A(B[1]), .B(n6460), .OUT(n6459) );
  NAND2 \gt_48/ULTI1_1  ( .A(\gt_48/AEQB [1]), .B(\gt_48/LTV [1]), .OUT(
        \gt_48/LTV2 [1]) );
  NAND2 \gt_48/ULTI2_1  ( .A(\gt_48/LTV1 [1]), .B(\gt_48/LTV2 [1]), .OUT(
        \gt_48/LTV [2]) );
  NOR2 \gt_48/ULTI0_2  ( .A(B[2]), .B(n6458), .OUT(n6457) );
  NAND2 \gt_48/ULTI1_2  ( .A(\gt_48/AEQB [2]), .B(\gt_48/LTV [2]), .OUT(
        \gt_48/LTV2 [2]) );
  NAND2 \gt_48/ULTI2_2  ( .A(\gt_48/LTV1 [2]), .B(\gt_48/LTV2 [2]), .OUT(
        \gt_48/LTV [3]) );
  NOR2 \gt_48/ULTI0_3  ( .A(B[3]), .B(n6456), .OUT(n6455) );
  NAND2 \gt_48/ULTI1_3  ( .A(\gt_48/AEQB [3]), .B(\gt_48/LTV [3]), .OUT(
        \gt_48/LTV2 [3]) );
  NAND2 \gt_48/ULTI2_3  ( .A(\gt_48/LTV1 [3]), .B(\gt_48/LTV2 [3]), .OUT(
        \gt_48/LTV [4]) );
  NOR2 \gt_48/ULTI0_4  ( .A(B[4]), .B(n6454), .OUT(n6453) );
  NAND2 \gt_48/ULTI1_4  ( .A(\gt_48/AEQB [4]), .B(\gt_48/LTV [4]), .OUT(
        \gt_48/LTV2 [4]) );
  NAND2 \gt_48/ULTI2_4  ( .A(\gt_48/LTV1 [4]), .B(\gt_48/LTV2 [4]), .OUT(
        \gt_48/LTV [5]) );
  NOR2 \gt_48/ULTI0_5  ( .A(B[5]), .B(n6452), .OUT(n6451) );
  NAND2 \gt_48/ULTI1_5  ( .A(\gt_48/AEQB [5]), .B(\gt_48/LTV [5]), .OUT(
        \gt_48/LTV2 [5]) );
  NAND2 \gt_48/ULTI2_5  ( .A(\gt_48/LTV1 [5]), .B(\gt_48/LTV2 [5]), .OUT(
        \gt_48/LTV [6]) );
  NOR2 \gt_48/ULTI0_6  ( .A(B[6]), .B(n6450), .OUT(n6449) );
  NAND2 \gt_48/ULTI1_6  ( .A(\gt_48/AEQB [6]), .B(\gt_48/LTV [6]), .OUT(
        \gt_48/LTV2 [6]) );
  NAND2 \gt_48/ULTI2_6  ( .A(\gt_48/LTV1 [6]), .B(\gt_48/LTV2 [6]), .OUT(
        \gt_48/LTV [7]) );
  NOR2 \gt_48/ULTI0_7  ( .A(B[7]), .B(n6448), .OUT(n6447) );
  NAND2 \gt_48/ULTI1_7  ( .A(\gt_48/AEQB [7]), .B(\gt_48/LTV [7]), .OUT(
        \gt_48/LTV2 [7]) );
  NAND2 \gt_48/ULTI2_7  ( .A(\gt_48/LTV1 [7]), .B(\gt_48/LTV2 [7]), .OUT(
        \gt_48/LTV [8]) );
  NOR2 \gt_48/ULTI0_8  ( .A(B[8]), .B(n6446), .OUT(n6445) );
  NAND2 \gt_48/ULTI1_8  ( .A(\gt_48/AEQB [8]), .B(\gt_48/LTV [8]), .OUT(
        \gt_48/LTV2 [8]) );
  NAND2 \gt_48/ULTI2_8  ( .A(\gt_48/LTV1 [8]), .B(\gt_48/LTV2 [8]), .OUT(
        \gt_48/LTV [9]) );
  NOR2 \gt_48/ULTI0_9  ( .A(B[9]), .B(n6444), .OUT(n6443) );
  NAND2 \gt_48/ULTI1_9  ( .A(\gt_48/AEQB [9]), .B(\gt_48/LTV [9]), .OUT(
        \gt_48/LTV2 [9]) );
  NAND2 \gt_48/ULTI2_9  ( .A(\gt_48/LTV1 [9]), .B(\gt_48/LTV2 [9]), .OUT(
        \gt_48/LTV [10]) );
  NOR2 \gt_48/ULTI0_10  ( .A(B[10]), .B(n6442), .OUT(n6441) );
  NAND2 \gt_48/ULTI1_10  ( .A(\gt_48/AEQB [10]), .B(\gt_48/LTV [10]), .OUT(
        \gt_48/LTV2 [10]) );
  NAND2 \gt_48/ULTI2_10  ( .A(\gt_48/LTV1 [10]), .B(\gt_48/LTV2 [10]), .OUT(
        \gt_48/LTV [11]) );
  NOR2 \gt_48/ULTI0_11  ( .A(B[11]), .B(n6440), .OUT(n6439) );
  NAND2 \gt_48/ULTI1_11  ( .A(\gt_48/AEQB [11]), .B(\gt_48/LTV [11]), .OUT(
        \gt_48/LTV2 [11]) );
  NAND2 \gt_48/ULTI2_11  ( .A(\gt_48/LTV1 [11]), .B(\gt_48/LTV2 [11]), .OUT(
        \gt_48/LTV [12]) );
  NOR2 \gt_48/ULTI0_12  ( .A(B[12]), .B(n6438), .OUT(n6437) );
  NAND2 \gt_48/ULTI1_12  ( .A(\gt_48/AEQB [12]), .B(\gt_48/LTV [12]), .OUT(
        \gt_48/LTV2 [12]) );
  NAND2 \gt_48/ULTI2_12  ( .A(\gt_48/LTV1 [12]), .B(\gt_48/LTV2 [12]), .OUT(
        \gt_48/LTV [13]) );
  NOR2 \gt_48/ULTI0_13  ( .A(B[13]), .B(n6436), .OUT(n6435) );
  NAND2 \gt_48/ULTI1_13  ( .A(\gt_48/AEQB [13]), .B(\gt_48/LTV [13]), .OUT(
        \gt_48/LTV2 [13]) );
  NAND2 \gt_48/ULTI2_13  ( .A(\gt_48/LTV1 [13]), .B(\gt_48/LTV2 [13]), .OUT(
        \gt_48/LTV [14]) );
  NOR2 \gt_48/ULTI0_14  ( .A(B[14]), .B(n6434), .OUT(n6433) );
  NAND2 \gt_48/ULTI1_14  ( .A(\gt_48/AEQB [14]), .B(\gt_48/LTV [14]), .OUT(
        \gt_48/LTV2 [14]) );
  NAND2 \gt_48/ULTI2_14  ( .A(\gt_48/LTV1 [14]), .B(\gt_48/LTV2 [14]), .OUT(
        \gt_48/LTV [15]) );
  NOR2 \gt_48/ULTI0_15  ( .A(B[15]), .B(n6432), .OUT(n6431) );
  NAND2 \gt_48/ULTI1_15  ( .A(\gt_48/AEQB [15]), .B(\gt_48/LTV [15]), .OUT(
        \gt_48/LTV2 [15]) );
  NAND2 \gt_48/ULTI2_15  ( .A(\gt_48/LTV1 [15]), .B(\gt_48/LTV2 [15]), .OUT(
        \gt_48/LTV [16]) );
  NOR2 \gt_48/ULTI0_16  ( .A(B[16]), .B(n6430), .OUT(n6429) );
  NAND2 \gt_48/ULTI1_16  ( .A(\gt_48/AEQB [16]), .B(\gt_48/LTV [16]), .OUT(
        \gt_48/LTV2 [16]) );
  NAND2 \gt_48/ULTI2_16  ( .A(\gt_48/LTV1 [16]), .B(\gt_48/LTV2 [16]), .OUT(
        \gt_48/LTV [17]) );
  NOR2 \gt_48/ULTI0_17  ( .A(B[17]), .B(n6428), .OUT(n6427) );
  NAND2 \gt_48/ULTI1_17  ( .A(\gt_48/AEQB [17]), .B(\gt_48/LTV [17]), .OUT(
        \gt_48/LTV2 [17]) );
  NAND2 \gt_48/ULTI2_17  ( .A(\gt_48/LTV1 [17]), .B(\gt_48/LTV2 [17]), .OUT(
        \gt_48/LTV [18]) );
  NOR2 \gt_48/ULTI0_18  ( .A(B[18]), .B(n6426), .OUT(n6425) );
  NAND2 \gt_48/ULTI1_18  ( .A(\gt_48/AEQB [18]), .B(\gt_48/LTV [18]), .OUT(
        \gt_48/LTV2 [18]) );
  NAND2 \gt_48/ULTI2_18  ( .A(\gt_48/LTV1 [18]), .B(\gt_48/LTV2 [18]), .OUT(
        \gt_48/LTV [19]) );
  NOR2 \gt_48/ULTI0_19  ( .A(B[19]), .B(n6424), .OUT(n6423) );
  NAND2 \gt_48/ULTI1_19  ( .A(\gt_48/AEQB [19]), .B(\gt_48/LTV [19]), .OUT(
        \gt_48/LTV2 [19]) );
  NAND2 \gt_48/ULTI2_19  ( .A(\gt_48/LTV1 [19]), .B(\gt_48/LTV2 [19]), .OUT(
        \gt_48/LTV [20]) );
  NOR2 \gt_48/ULTI0_20  ( .A(B[20]), .B(n6422), .OUT(n6421) );
  NAND2 \gt_48/ULTI1_20  ( .A(\gt_48/AEQB [20]), .B(\gt_48/LTV [20]), .OUT(
        \gt_48/LTV2 [20]) );
  NAND2 \gt_48/ULTI2_20  ( .A(\gt_48/LTV1 [20]), .B(\gt_48/LTV2 [20]), .OUT(
        \gt_48/LTV [21]) );
  NOR2 \gt_48/ULTI0_21  ( .A(B[21]), .B(n6420), .OUT(n6419) );
  NAND2 \gt_48/ULTI1_21  ( .A(\gt_48/AEQB [21]), .B(\gt_48/LTV [21]), .OUT(
        \gt_48/LTV2 [21]) );
  NAND2 \gt_48/ULTI2_21  ( .A(\gt_48/LTV1 [21]), .B(\gt_48/LTV2 [21]), .OUT(
        \gt_48/LTV [22]) );
  NOR2 \gt_48/ULTI0_22  ( .A(B[22]), .B(n6418), .OUT(n6417) );
  NAND2 \gt_48/ULTI1_22  ( .A(\gt_48/AEQB [22]), .B(\gt_48/LTV [22]), .OUT(
        \gt_48/LTV2 [22]) );
  NAND2 \gt_48/ULTI2_22  ( .A(\gt_48/LTV1 [22]), .B(\gt_48/LTV2 [22]), .OUT(
        \gt_48/LTV [23]) );
  NOR2 \gt_48/ULTI0_23  ( .A(B[23]), .B(n6416), .OUT(n6415) );
  NAND2 \gt_48/ULTI1_23  ( .A(\gt_48/AEQB [23]), .B(\gt_48/LTV [23]), .OUT(
        \gt_48/LTV2 [23]) );
  NAND2 \gt_48/ULTI2_23  ( .A(\gt_48/LTV1 [23]), .B(\gt_48/LTV2 [23]), .OUT(
        \gt_48/LTV [24]) );
  NOR2 \gt_48/ULTI0_24  ( .A(B[24]), .B(n6414), .OUT(n6413) );
  NAND2 \gt_48/ULTI1_24  ( .A(\gt_48/AEQB [24]), .B(\gt_48/LTV [24]), .OUT(
        \gt_48/LTV2 [24]) );
  NAND2 \gt_48/ULTI2_24  ( .A(\gt_48/LTV1 [24]), .B(\gt_48/LTV2 [24]), .OUT(
        \gt_48/LTV [25]) );
  NOR2 \gt_48/ULTI0_25  ( .A(B[25]), .B(n6412), .OUT(n6411) );
  NAND2 \gt_48/ULTI1_25  ( .A(\gt_48/AEQB [25]), .B(\gt_48/LTV [25]), .OUT(
        \gt_48/LTV2 [25]) );
  NAND2 \gt_48/ULTI2_25  ( .A(\gt_48/LTV1 [25]), .B(\gt_48/LTV2 [25]), .OUT(
        \gt_48/LTV [26]) );
  NOR2 \gt_48/ULTI0_26  ( .A(B[26]), .B(n6410), .OUT(n6409) );
  NAND2 \gt_48/ULTI1_26  ( .A(\gt_48/AEQB [26]), .B(\gt_48/LTV [26]), .OUT(
        \gt_48/LTV2 [26]) );
  NAND2 \gt_48/ULTI2_26  ( .A(\gt_48/LTV1 [26]), .B(\gt_48/LTV2 [26]), .OUT(
        \gt_48/LTV [27]) );
  NOR2 \gt_48/ULTI0_27  ( .A(B[27]), .B(n6408), .OUT(n6407) );
  NAND2 \gt_48/ULTI1_27  ( .A(\gt_48/AEQB [27]), .B(\gt_48/LTV [27]), .OUT(
        \gt_48/LTV2 [27]) );
  NAND2 \gt_48/ULTI2_27  ( .A(\gt_48/LTV1 [27]), .B(\gt_48/LTV2 [27]), .OUT(
        \gt_48/LTV [28]) );
  NOR2 \gt_48/ULTI0_28  ( .A(B[28]), .B(n6406), .OUT(n6405) );
  NAND2 \gt_48/ULTI1_28  ( .A(\gt_48/AEQB [28]), .B(\gt_48/LTV [28]), .OUT(
        \gt_48/LTV2 [28]) );
  NAND2 \gt_48/ULTI2_28  ( .A(\gt_48/LTV1 [28]), .B(\gt_48/LTV2 [28]), .OUT(
        \gt_48/LTV [29]) );
  NOR2 \gt_48/ULTI0_29  ( .A(B[29]), .B(n6404), .OUT(n6403) );
  NAND2 \gt_48/ULTI1_29  ( .A(\gt_48/AEQB [29]), .B(\gt_48/LTV [29]), .OUT(
        \gt_48/LTV2 [29]) );
  NAND2 \gt_48/ULTI2_29  ( .A(\gt_48/LTV1 [29]), .B(\gt_48/LTV2 [29]), .OUT(
        \gt_48/LTV [30]) );
  NOR2 \gt_48/ULTI0_30  ( .A(B[30]), .B(n6402), .OUT(n6401) );
  NAND2 \gt_48/ULTI1_30  ( .A(\gt_48/AEQB [30]), .B(\gt_48/LTV [30]), .OUT(
        \gt_48/LTV2 [30]) );
  NAND2 \gt_48/ULTI2_30  ( .A(\gt_48/LTV1 [30]), .B(\gt_48/LTV2 [30]), .OUT(
        \gt_48/LTV [31]) );
  NOR2 \gt_48/ULTI0  ( .A(\gt_48/SA ), .B(n6400), .OUT(n6399) );
  NAND2 \gt_48/ULTI1  ( .A(\gt_48/AEQB [31]), .B(\gt_48/LTV [31]), .OUT(
        \gt_48/LTV2 [31]) );
  NAND2 \gt_48/ULTI2  ( .A(\gt_48/LTV1 [31]), .B(\gt_48/LTV2 [31]), .OUT(N221)
         );
  INV U316 ( .IN(\gt_48/LTV1 [0]), .OUT(\gt_48/LTV [1]) );
  INV U317 ( .IN(\mult_49/A1[0] ), .OUT(n6463) );
  INV U318 ( .IN(\mult_49/A1[1] ), .OUT(n6464) );
  INV U319 ( .IN(n6463), .OUT(N224) );
  INV U320 ( .IN(\mult_49/A1[2] ), .OUT(n6465) );
  INV U321 ( .IN(n6464), .OUT(N225) );
  INV U322 ( .IN(\mult_49/A1[3] ), .OUT(n6466) );
  INV U323 ( .IN(n6465), .OUT(N226) );
  INV U324 ( .IN(\mult_49/A1[4] ), .OUT(n6467) );
  INV U325 ( .IN(n6466), .OUT(N227) );
  INV U326 ( .IN(\mult_49/A1[5] ), .OUT(n6468) );
  INV U327 ( .IN(n6467), .OUT(N228) );
  INV U328 ( .IN(\mult_49/A1[6] ), .OUT(n6469) );
  INV U329 ( .IN(n6468), .OUT(N229) );
  INV U330 ( .IN(\mult_49/A1[7] ), .OUT(n6470) );
  INV U331 ( .IN(n6469), .OUT(N230) );
  INV U332 ( .IN(\mult_49/A1[8] ), .OUT(n6471) );
  INV U333 ( .IN(n6470), .OUT(N231) );
  INV U334 ( .IN(\mult_49/A1[9] ), .OUT(n6472) );
  INV U335 ( .IN(n6471), .OUT(N232) );
  INV U336 ( .IN(\mult_49/A1[10] ), .OUT(n6473) );
  INV U337 ( .IN(n6472), .OUT(N233) );
  INV U338 ( .IN(\mult_49/A1[11] ), .OUT(n6474) );
  INV U339 ( .IN(n6473), .OUT(N234) );
  INV U340 ( .IN(\mult_49/A1[12] ), .OUT(n6475) );
  INV U341 ( .IN(n6474), .OUT(N235) );
  INV U342 ( .IN(\mult_49/A1[13] ), .OUT(n6476) );
  INV U343 ( .IN(n6475), .OUT(N236) );
  INV U344 ( .IN(\mult_49/A1[14] ), .OUT(n6477) );
  INV U345 ( .IN(n6476), .OUT(N237) );
  INV U346 ( .IN(\mult_49/A1[15] ), .OUT(n6478) );
  INV U347 ( .IN(n6477), .OUT(N238) );
  INV U348 ( .IN(\mult_49/A1[16] ), .OUT(n6479) );
  INV U349 ( .IN(n6478), .OUT(N239) );
  INV U350 ( .IN(\mult_49/A1[17] ), .OUT(n6480) );
  INV U351 ( .IN(n6479), .OUT(N240) );
  INV U352 ( .IN(\mult_49/A1[18] ), .OUT(n6481) );
  INV U353 ( .IN(n6480), .OUT(N241) );
  INV U354 ( .IN(\mult_49/A1[19] ), .OUT(n6482) );
  INV U355 ( .IN(n6481), .OUT(N242) );
  INV U356 ( .IN(\mult_49/A1[20] ), .OUT(n6483) );
  INV U357 ( .IN(n6482), .OUT(N243) );
  INV U358 ( .IN(\mult_49/A1[21] ), .OUT(n6484) );
  INV U359 ( .IN(n6483), .OUT(N244) );
  INV U360 ( .IN(\mult_49/A1[22] ), .OUT(n6485) );
  INV U361 ( .IN(n6484), .OUT(N245) );
  INV U362 ( .IN(\mult_49/A1[23] ), .OUT(n6486) );
  INV U363 ( .IN(n6485), .OUT(N246) );
  INV U364 ( .IN(\mult_49/A1[24] ), .OUT(n6487) );
  INV U365 ( .IN(n6486), .OUT(N247) );
  INV U366 ( .IN(\mult_49/A1[25] ), .OUT(n6488) );
  INV U367 ( .IN(n6487), .OUT(N248) );
  INV U368 ( .IN(\mult_49/A1[26] ), .OUT(n6489) );
  INV U369 ( .IN(n6488), .OUT(N249) );
  INV U370 ( .IN(\mult_49/A1[27] ), .OUT(n6490) );
  INV U371 ( .IN(n6489), .OUT(N250) );
  INV U372 ( .IN(\mult_49/A1[28] ), .OUT(n6491) );
  INV U373 ( .IN(n6490), .OUT(N251) );
  INV U374 ( .IN(\mult_49/A1[29] ), .OUT(n6492) );
  INV U375 ( .IN(n6491), .OUT(N252) );
  INV U376 ( .IN(n6492), .OUT(N253) );
  NAND2 U377 ( .A(n289), .B(n290), .OUT(N93) );
  INV U378 ( .IN(B[0]), .OUT(\mult_49/B_notx[0] ) );
  INV U379 ( .IN(A[0]), .OUT(\mult_49/A_notx[0] ) );
  NOR2 U380 ( .A(n292), .B(n293), .OUT(n291) );
  INV U381 ( .IN(\mult_49/ab[2][9] ), .OUT(n294) );
  INV U382 ( .IN(\mult_49/ab[2][8] ), .OUT(n295) );
  NOR2 U383 ( .A(n297), .B(n298), .OUT(n296) );
  INV U384 ( .IN(\mult_49/ab[3][8] ), .OUT(n299) );
  NAND2 U385 ( .A(n301), .B(n302), .OUT(n300) );
  INV U386 ( .IN(\mult_49/ab[2][7] ), .OUT(n303) );
  NOR2 U387 ( .A(n305), .B(n306), .OUT(n304) );
  NAND2 U388 ( .A(n308), .B(n309), .OUT(n307) );
  INV U389 ( .IN(\mult_49/ab[3][7] ), .OUT(n310) );
  INV U390 ( .IN(\mult_49/ab[4][7] ), .OUT(n311) );
  NAND2 U391 ( .A(n313), .B(n314), .OUT(n312) );
  INV U392 ( .IN(\mult_49/ab[2][6] ), .OUT(n315) );
  NOR2 U393 ( .A(n317), .B(n318), .OUT(n316) );
  NAND2 U394 ( .A(n320), .B(n321), .OUT(n319) );
  INV U395 ( .IN(\mult_49/ab[3][6] ), .OUT(n322) );
  NAND2 U396 ( .A(n324), .B(n325), .OUT(n323) );
  INV U397 ( .IN(\mult_49/ab[4][6] ), .OUT(n326) );
  INV U398 ( .IN(\mult_49/ab[5][6] ), .OUT(n327) );
  NAND2 U399 ( .A(n329), .B(n330), .OUT(n328) );
  INV U400 ( .IN(\mult_49/ab[2][5] ), .OUT(n331) );
  NOR2 U401 ( .A(n333), .B(n334), .OUT(n332) );
  NAND2 U402 ( .A(n336), .B(n337), .OUT(n335) );
  INV U403 ( .IN(\mult_49/ab[3][5] ), .OUT(n338) );
  NAND2 U404 ( .A(n340), .B(n341), .OUT(n339) );
  INV U405 ( .IN(\mult_49/ab[4][5] ), .OUT(n342) );
  NAND2 U406 ( .A(n344), .B(n345), .OUT(n343) );
  INV U407 ( .IN(\mult_49/ab[5][5] ), .OUT(n346) );
  INV U408 ( .IN(\mult_49/ab[6][5] ), .OUT(n347) );
  NAND2 U409 ( .A(n349), .B(n350), .OUT(n348) );
  INV U410 ( .IN(\mult_49/ab[2][4] ), .OUT(n351) );
  NOR2 U411 ( .A(n353), .B(n354), .OUT(n352) );
  NAND2 U412 ( .A(n356), .B(n357), .OUT(n355) );
  INV U413 ( .IN(\mult_49/ab[3][4] ), .OUT(n358) );
  NAND2 U414 ( .A(n360), .B(n361), .OUT(n359) );
  INV U415 ( .IN(\mult_49/ab[4][4] ), .OUT(n362) );
  NAND2 U416 ( .A(n364), .B(n365), .OUT(n363) );
  INV U417 ( .IN(\mult_49/ab[5][4] ), .OUT(n366) );
  NAND2 U418 ( .A(n368), .B(n369), .OUT(n367) );
  INV U419 ( .IN(\mult_49/ab[6][4] ), .OUT(n370) );
  INV U420 ( .IN(\mult_49/ab[7][4] ), .OUT(n371) );
  NAND2 U421 ( .A(n373), .B(n374), .OUT(n372) );
  INV U422 ( .IN(\mult_49/ab[2][3] ), .OUT(n375) );
  NOR2 U423 ( .A(n377), .B(n378), .OUT(n376) );
  NAND2 U424 ( .A(n380), .B(n381), .OUT(n379) );
  INV U425 ( .IN(\mult_49/ab[3][3] ), .OUT(n382) );
  NAND2 U426 ( .A(n384), .B(n385), .OUT(n383) );
  INV U427 ( .IN(\mult_49/ab[4][3] ), .OUT(n386) );
  NAND2 U428 ( .A(n388), .B(n389), .OUT(n387) );
  INV U429 ( .IN(\mult_49/ab[5][3] ), .OUT(n390) );
  NAND2 U430 ( .A(n392), .B(n393), .OUT(n391) );
  INV U431 ( .IN(\mult_49/ab[6][3] ), .OUT(n394) );
  NAND2 U432 ( .A(n396), .B(n397), .OUT(n395) );
  INV U433 ( .IN(\mult_49/ab[7][3] ), .OUT(n398) );
  INV U434 ( .IN(\mult_49/ab[8][3] ), .OUT(n399) );
  NAND2 U435 ( .A(n401), .B(n402), .OUT(n400) );
  INV U436 ( .IN(\mult_49/ab[2][2] ), .OUT(n403) );
  NOR2 U437 ( .A(n405), .B(n406), .OUT(n404) );
  NAND2 U438 ( .A(n408), .B(n409), .OUT(n407) );
  INV U439 ( .IN(\mult_49/ab[3][2] ), .OUT(n410) );
  NAND2 U440 ( .A(n412), .B(n413), .OUT(n411) );
  INV U441 ( .IN(\mult_49/ab[4][2] ), .OUT(n414) );
  NAND2 U442 ( .A(n416), .B(n417), .OUT(n415) );
  INV U443 ( .IN(\mult_49/ab[5][2] ), .OUT(n418) );
  NAND2 U444 ( .A(n420), .B(n421), .OUT(n419) );
  INV U445 ( .IN(\mult_49/ab[6][2] ), .OUT(n422) );
  NAND2 U446 ( .A(n424), .B(n425), .OUT(n423) );
  INV U447 ( .IN(\mult_49/ab[7][2] ), .OUT(n426) );
  NAND2 U448 ( .A(n428), .B(n429), .OUT(n427) );
  INV U449 ( .IN(\mult_49/ab[8][2] ), .OUT(n430) );
  INV U450 ( .IN(\mult_49/ab[9][2] ), .OUT(n431) );
  NAND2 U451 ( .A(n433), .B(n434), .OUT(n432) );
  INV U452 ( .IN(\mult_49/ab[2][1] ), .OUT(n435) );
  NOR2 U453 ( .A(n437), .B(n438), .OUT(n436) );
  NAND2 U454 ( .A(n440), .B(n441), .OUT(n439) );
  INV U455 ( .IN(\mult_49/ab[3][1] ), .OUT(n442) );
  NAND2 U456 ( .A(n444), .B(n445), .OUT(n443) );
  INV U457 ( .IN(\mult_49/ab[4][1] ), .OUT(n446) );
  NAND2 U458 ( .A(n448), .B(n449), .OUT(n447) );
  INV U459 ( .IN(\mult_49/ab[5][1] ), .OUT(n450) );
  NAND2 U460 ( .A(n452), .B(n453), .OUT(n451) );
  INV U461 ( .IN(\mult_49/ab[6][1] ), .OUT(n454) );
  NAND2 U462 ( .A(n456), .B(n457), .OUT(n455) );
  INV U463 ( .IN(\mult_49/ab[7][1] ), .OUT(n458) );
  NAND2 U464 ( .A(n460), .B(n461), .OUT(n459) );
  INV U465 ( .IN(\mult_49/ab[8][1] ), .OUT(n462) );
  NAND2 U466 ( .A(n464), .B(n465), .OUT(n463) );
  INV U467 ( .IN(\mult_49/ab[9][1] ), .OUT(n466) );
  INV U468 ( .IN(\mult_49/ab[10][1] ), .OUT(n467) );
  NAND2 U469 ( .A(n469), .B(n470), .OUT(n468) );
  INV U470 ( .IN(\mult_49/ab[2][0] ), .OUT(n471) );
  NOR2 U471 ( .A(n473), .B(n474), .OUT(n472) );
  NAND2 U472 ( .A(n476), .B(n477), .OUT(n475) );
  INV U473 ( .IN(\mult_49/ab[3][0] ), .OUT(n478) );
  NAND2 U474 ( .A(n480), .B(n481), .OUT(n479) );
  INV U475 ( .IN(\mult_49/ab[4][0] ), .OUT(n482) );
  NAND2 U476 ( .A(n484), .B(n485), .OUT(n483) );
  INV U477 ( .IN(\mult_49/ab[5][0] ), .OUT(n486) );
  NAND2 U478 ( .A(n488), .B(n489), .OUT(n487) );
  INV U479 ( .IN(\mult_49/ab[6][0] ), .OUT(n490) );
  NAND2 U480 ( .A(n492), .B(n493), .OUT(n491) );
  INV U481 ( .IN(\mult_49/ab[7][0] ), .OUT(n494) );
  NAND2 U482 ( .A(n496), .B(n497), .OUT(n495) );
  INV U483 ( .IN(\mult_49/ab[8][0] ), .OUT(n498) );
  NAND2 U484 ( .A(n500), .B(n501), .OUT(n499) );
  INV U485 ( .IN(\mult_49/ab[9][0] ), .OUT(n502) );
  NAND2 U486 ( .A(n504), .B(n505), .OUT(n503) );
  INV U487 ( .IN(\mult_49/ab[10][0] ), .OUT(n506) );
  INV U488 ( .IN(\mult_49/ab[11][0] ), .OUT(n507) );
  NAND2 U489 ( .A(n509), .B(n510), .OUT(n508) );
  NAND2 U490 ( .A(n512), .B(n513), .OUT(n511) );
  NOR2 U491 ( .A(n515), .B(n516), .OUT(n514) );
  INV U492 ( .IN(\mult_49/ab[2][10] ), .OUT(n517) );
  INV U493 ( .IN(\mult_49/ab[3][9] ), .OUT(n518) );
  NAND2 U494 ( .A(n520), .B(n521), .OUT(n519) );
  INV U495 ( .IN(\mult_49/ab[4][8] ), .OUT(n522) );
  NAND2 U496 ( .A(n524), .B(n525), .OUT(n523) );
  INV U497 ( .IN(\mult_49/ab[5][7] ), .OUT(n526) );
  NAND2 U498 ( .A(n528), .B(n529), .OUT(n527) );
  INV U499 ( .IN(\mult_49/ab[6][6] ), .OUT(n530) );
  NAND2 U500 ( .A(n532), .B(n533), .OUT(n531) );
  INV U501 ( .IN(\mult_49/ab[7][5] ), .OUT(n534) );
  NAND2 U502 ( .A(n536), .B(n537), .OUT(n535) );
  INV U503 ( .IN(\mult_49/ab[8][4] ), .OUT(n538) );
  NAND2 U504 ( .A(n540), .B(n541), .OUT(n539) );
  INV U505 ( .IN(\mult_49/ab[9][3] ), .OUT(n542) );
  NAND2 U506 ( .A(n544), .B(n545), .OUT(n543) );
  INV U507 ( .IN(\mult_49/ab[10][2] ), .OUT(n546) );
  NAND2 U508 ( .A(n548), .B(n549), .OUT(n547) );
  NOR2 U509 ( .A(n551), .B(n552), .OUT(n550) );
  INV U510 ( .IN(\mult_49/ab[2][11] ), .OUT(n553) );
  INV U511 ( .IN(\mult_49/ab[3][10] ), .OUT(n554) );
  NAND2 U512 ( .A(n556), .B(n557), .OUT(n555) );
  INV U513 ( .IN(\mult_49/ab[4][9] ), .OUT(n558) );
  NAND2 U514 ( .A(n560), .B(n561), .OUT(n559) );
  INV U515 ( .IN(\mult_49/ab[5][8] ), .OUT(n562) );
  NAND2 U516 ( .A(n564), .B(n565), .OUT(n563) );
  INV U517 ( .IN(\mult_49/ab[6][7] ), .OUT(n566) );
  NAND2 U518 ( .A(n568), .B(n569), .OUT(n567) );
  INV U519 ( .IN(\mult_49/ab[7][6] ), .OUT(n570) );
  NAND2 U520 ( .A(n572), .B(n573), .OUT(n571) );
  INV U521 ( .IN(\mult_49/ab[8][5] ), .OUT(n574) );
  NAND2 U522 ( .A(n576), .B(n577), .OUT(n575) );
  INV U523 ( .IN(\mult_49/ab[9][4] ), .OUT(n578) );
  NAND2 U524 ( .A(n580), .B(n581), .OUT(n579) );
  INV U525 ( .IN(\mult_49/ab[10][3] ), .OUT(n582) );
  NAND2 U526 ( .A(n584), .B(n585), .OUT(n583) );
  INV U527 ( .IN(\mult_49/ab[11][2] ), .OUT(n586) );
  NAND2 U528 ( .A(n588), .B(n589), .OUT(n587) );
  NOR2 U529 ( .A(n591), .B(n592), .OUT(n590) );
  INV U530 ( .IN(\mult_49/ab[2][12] ), .OUT(n593) );
  INV U531 ( .IN(\mult_49/ab[3][11] ), .OUT(n594) );
  NAND2 U532 ( .A(n596), .B(n597), .OUT(n595) );
  INV U533 ( .IN(\mult_49/ab[4][10] ), .OUT(n598) );
  NAND2 U534 ( .A(n600), .B(n601), .OUT(n599) );
  INV U535 ( .IN(\mult_49/ab[5][9] ), .OUT(n602) );
  NAND2 U536 ( .A(n604), .B(n605), .OUT(n603) );
  INV U537 ( .IN(\mult_49/ab[6][8] ), .OUT(n606) );
  NAND2 U538 ( .A(n608), .B(n609), .OUT(n607) );
  INV U539 ( .IN(\mult_49/ab[7][7] ), .OUT(n610) );
  NAND2 U540 ( .A(n612), .B(n613), .OUT(n611) );
  INV U541 ( .IN(\mult_49/ab[8][6] ), .OUT(n614) );
  NAND2 U542 ( .A(n616), .B(n617), .OUT(n615) );
  INV U543 ( .IN(\mult_49/ab[9][5] ), .OUT(n618) );
  NAND2 U544 ( .A(n620), .B(n621), .OUT(n619) );
  INV U545 ( .IN(\mult_49/ab[10][4] ), .OUT(n622) );
  NAND2 U546 ( .A(n624), .B(n625), .OUT(n623) );
  INV U547 ( .IN(\mult_49/ab[11][3] ), .OUT(n626) );
  NAND2 U548 ( .A(n628), .B(n629), .OUT(n627) );
  INV U549 ( .IN(\mult_49/ab[12][2] ), .OUT(n630) );
  NAND2 U550 ( .A(n632), .B(n633), .OUT(n631) );
  NOR2 U551 ( .A(n635), .B(n636), .OUT(n634) );
  INV U552 ( .IN(\mult_49/ab[2][13] ), .OUT(n637) );
  INV U553 ( .IN(\mult_49/ab[3][12] ), .OUT(n638) );
  NAND2 U554 ( .A(n640), .B(n641), .OUT(n639) );
  INV U555 ( .IN(\mult_49/ab[4][11] ), .OUT(n642) );
  NAND2 U556 ( .A(n644), .B(n645), .OUT(n643) );
  INV U557 ( .IN(\mult_49/ab[5][10] ), .OUT(n646) );
  NAND2 U558 ( .A(n648), .B(n649), .OUT(n647) );
  INV U559 ( .IN(\mult_49/ab[6][9] ), .OUT(n650) );
  NAND2 U560 ( .A(n652), .B(n653), .OUT(n651) );
  INV U561 ( .IN(\mult_49/ab[7][8] ), .OUT(n654) );
  NAND2 U562 ( .A(n656), .B(n657), .OUT(n655) );
  INV U563 ( .IN(\mult_49/ab[8][7] ), .OUT(n658) );
  NAND2 U564 ( .A(n660), .B(n661), .OUT(n659) );
  INV U565 ( .IN(\mult_49/ab[9][6] ), .OUT(n662) );
  NAND2 U566 ( .A(n664), .B(n665), .OUT(n663) );
  INV U567 ( .IN(\mult_49/ab[10][5] ), .OUT(n666) );
  NAND2 U568 ( .A(n668), .B(n669), .OUT(n667) );
  INV U569 ( .IN(\mult_49/ab[11][4] ), .OUT(n670) );
  NAND2 U570 ( .A(n672), .B(n673), .OUT(n671) );
  INV U571 ( .IN(\mult_49/ab[12][3] ), .OUT(n674) );
  NAND2 U572 ( .A(n676), .B(n677), .OUT(n675) );
  INV U573 ( .IN(\mult_49/ab[13][2] ), .OUT(n678) );
  NAND2 U574 ( .A(n680), .B(n681), .OUT(n679) );
  NOR2 U575 ( .A(n683), .B(n684), .OUT(n682) );
  INV U576 ( .IN(\mult_49/ab[2][14] ), .OUT(n685) );
  INV U577 ( .IN(\mult_49/ab[3][13] ), .OUT(n686) );
  NAND2 U578 ( .A(n688), .B(n689), .OUT(n687) );
  INV U579 ( .IN(\mult_49/ab[4][12] ), .OUT(n690) );
  NAND2 U580 ( .A(n692), .B(n693), .OUT(n691) );
  INV U581 ( .IN(\mult_49/ab[5][11] ), .OUT(n694) );
  NAND2 U582 ( .A(n696), .B(n697), .OUT(n695) );
  INV U583 ( .IN(\mult_49/ab[6][10] ), .OUT(n698) );
  NAND2 U584 ( .A(n700), .B(n701), .OUT(n699) );
  INV U585 ( .IN(\mult_49/ab[7][9] ), .OUT(n702) );
  NAND2 U586 ( .A(n704), .B(n705), .OUT(n703) );
  INV U587 ( .IN(\mult_49/ab[8][8] ), .OUT(n706) );
  NAND2 U588 ( .A(n708), .B(n709), .OUT(n707) );
  INV U589 ( .IN(\mult_49/ab[9][7] ), .OUT(n710) );
  NAND2 U590 ( .A(n712), .B(n713), .OUT(n711) );
  INV U591 ( .IN(\mult_49/ab[10][6] ), .OUT(n714) );
  NAND2 U592 ( .A(n716), .B(n717), .OUT(n715) );
  INV U593 ( .IN(\mult_49/ab[11][5] ), .OUT(n718) );
  NAND2 U594 ( .A(n720), .B(n721), .OUT(n719) );
  INV U595 ( .IN(\mult_49/ab[12][4] ), .OUT(n722) );
  NAND2 U596 ( .A(n724), .B(n725), .OUT(n723) );
  INV U597 ( .IN(\mult_49/ab[13][3] ), .OUT(n726) );
  NAND2 U598 ( .A(n728), .B(n729), .OUT(n727) );
  INV U599 ( .IN(\mult_49/ab[14][2] ), .OUT(n730) );
  NAND2 U600 ( .A(n732), .B(n733), .OUT(n731) );
  NOR2 U601 ( .A(n735), .B(n736), .OUT(n734) );
  INV U602 ( .IN(\mult_49/ab[2][15] ), .OUT(n737) );
  INV U603 ( .IN(\mult_49/ab[3][14] ), .OUT(n738) );
  NAND2 U604 ( .A(n740), .B(n741), .OUT(n739) );
  INV U605 ( .IN(\mult_49/ab[4][13] ), .OUT(n742) );
  NAND2 U606 ( .A(n744), .B(n745), .OUT(n743) );
  INV U607 ( .IN(\mult_49/ab[5][12] ), .OUT(n746) );
  NAND2 U608 ( .A(n748), .B(n749), .OUT(n747) );
  INV U609 ( .IN(\mult_49/ab[6][11] ), .OUT(n750) );
  NAND2 U610 ( .A(n752), .B(n753), .OUT(n751) );
  INV U611 ( .IN(\mult_49/ab[7][10] ), .OUT(n754) );
  NAND2 U612 ( .A(n756), .B(n757), .OUT(n755) );
  INV U613 ( .IN(\mult_49/ab[8][9] ), .OUT(n758) );
  NAND2 U614 ( .A(n760), .B(n761), .OUT(n759) );
  INV U615 ( .IN(\mult_49/ab[9][8] ), .OUT(n762) );
  NAND2 U616 ( .A(n764), .B(n765), .OUT(n763) );
  INV U617 ( .IN(\mult_49/ab[10][7] ), .OUT(n766) );
  NAND2 U618 ( .A(n768), .B(n769), .OUT(n767) );
  INV U619 ( .IN(\mult_49/ab[11][6] ), .OUT(n770) );
  NAND2 U620 ( .A(n772), .B(n773), .OUT(n771) );
  INV U621 ( .IN(\mult_49/ab[12][5] ), .OUT(n774) );
  NAND2 U622 ( .A(n776), .B(n777), .OUT(n775) );
  INV U623 ( .IN(\mult_49/ab[13][4] ), .OUT(n778) );
  NAND2 U624 ( .A(n780), .B(n781), .OUT(n779) );
  INV U625 ( .IN(\mult_49/ab[14][3] ), .OUT(n782) );
  NAND2 U626 ( .A(n784), .B(n785), .OUT(n783) );
  INV U627 ( .IN(\mult_49/ab[15][2] ), .OUT(n786) );
  NAND2 U628 ( .A(n788), .B(n789), .OUT(n787) );
  NOR2 U629 ( .A(n791), .B(n792), .OUT(n790) );
  INV U630 ( .IN(\mult_49/ab[2][16] ), .OUT(n793) );
  INV U631 ( .IN(\mult_49/ab[3][15] ), .OUT(n794) );
  NAND2 U632 ( .A(n796), .B(n797), .OUT(n795) );
  INV U633 ( .IN(\mult_49/ab[4][14] ), .OUT(n798) );
  NAND2 U634 ( .A(n800), .B(n801), .OUT(n799) );
  INV U635 ( .IN(\mult_49/ab[5][13] ), .OUT(n802) );
  NAND2 U636 ( .A(n804), .B(n805), .OUT(n803) );
  INV U637 ( .IN(\mult_49/ab[6][12] ), .OUT(n806) );
  NAND2 U638 ( .A(n808), .B(n809), .OUT(n807) );
  INV U639 ( .IN(\mult_49/ab[7][11] ), .OUT(n810) );
  NAND2 U640 ( .A(n812), .B(n813), .OUT(n811) );
  INV U641 ( .IN(\mult_49/ab[8][10] ), .OUT(n814) );
  NAND2 U642 ( .A(n816), .B(n817), .OUT(n815) );
  INV U643 ( .IN(\mult_49/ab[9][9] ), .OUT(n818) );
  NAND2 U644 ( .A(n820), .B(n821), .OUT(n819) );
  INV U645 ( .IN(\mult_49/ab[10][8] ), .OUT(n822) );
  NAND2 U646 ( .A(n824), .B(n825), .OUT(n823) );
  INV U647 ( .IN(\mult_49/ab[11][7] ), .OUT(n826) );
  NAND2 U648 ( .A(n828), .B(n829), .OUT(n827) );
  INV U649 ( .IN(\mult_49/ab[12][6] ), .OUT(n830) );
  NAND2 U650 ( .A(n832), .B(n833), .OUT(n831) );
  INV U651 ( .IN(\mult_49/ab[13][5] ), .OUT(n834) );
  NAND2 U652 ( .A(n836), .B(n837), .OUT(n835) );
  INV U653 ( .IN(\mult_49/ab[14][4] ), .OUT(n838) );
  NAND2 U654 ( .A(n840), .B(n841), .OUT(n839) );
  INV U655 ( .IN(\mult_49/ab[15][3] ), .OUT(n842) );
  NAND2 U656 ( .A(n844), .B(n845), .OUT(n843) );
  INV U657 ( .IN(\mult_49/ab[16][2] ), .OUT(n846) );
  NAND2 U658 ( .A(n848), .B(n849), .OUT(n847) );
  NOR2 U659 ( .A(n851), .B(n852), .OUT(n850) );
  INV U660 ( .IN(\mult_49/ab[2][17] ), .OUT(n853) );
  INV U661 ( .IN(\mult_49/ab[3][16] ), .OUT(n854) );
  NAND2 U662 ( .A(n856), .B(n857), .OUT(n855) );
  INV U663 ( .IN(\mult_49/ab[4][15] ), .OUT(n858) );
  NAND2 U664 ( .A(n860), .B(n861), .OUT(n859) );
  INV U665 ( .IN(\mult_49/ab[5][14] ), .OUT(n862) );
  NAND2 U666 ( .A(n864), .B(n865), .OUT(n863) );
  INV U667 ( .IN(\mult_49/ab[6][13] ), .OUT(n866) );
  NAND2 U668 ( .A(n868), .B(n869), .OUT(n867) );
  INV U669 ( .IN(\mult_49/ab[7][12] ), .OUT(n870) );
  NAND2 U670 ( .A(n872), .B(n873), .OUT(n871) );
  INV U671 ( .IN(\mult_49/ab[8][11] ), .OUT(n874) );
  NAND2 U672 ( .A(n876), .B(n877), .OUT(n875) );
  INV U673 ( .IN(\mult_49/ab[9][10] ), .OUT(n878) );
  NAND2 U674 ( .A(n880), .B(n881), .OUT(n879) );
  INV U675 ( .IN(\mult_49/ab[10][9] ), .OUT(n882) );
  NAND2 U676 ( .A(n884), .B(n885), .OUT(n883) );
  INV U677 ( .IN(\mult_49/ab[11][8] ), .OUT(n886) );
  NAND2 U678 ( .A(n888), .B(n889), .OUT(n887) );
  INV U679 ( .IN(\mult_49/ab[12][7] ), .OUT(n890) );
  NAND2 U680 ( .A(n892), .B(n893), .OUT(n891) );
  INV U681 ( .IN(\mult_49/ab[13][6] ), .OUT(n894) );
  NAND2 U682 ( .A(n896), .B(n897), .OUT(n895) );
  INV U683 ( .IN(\mult_49/ab[14][5] ), .OUT(n898) );
  NAND2 U684 ( .A(n900), .B(n901), .OUT(n899) );
  INV U685 ( .IN(\mult_49/ab[15][4] ), .OUT(n902) );
  NAND2 U686 ( .A(n904), .B(n905), .OUT(n903) );
  INV U687 ( .IN(\mult_49/ab[16][3] ), .OUT(n906) );
  NAND2 U688 ( .A(n908), .B(n909), .OUT(n907) );
  INV U689 ( .IN(\mult_49/ab[17][2] ), .OUT(n910) );
  NAND2 U690 ( .A(n912), .B(n913), .OUT(n911) );
  NOR2 U691 ( .A(n915), .B(n916), .OUT(n914) );
  INV U692 ( .IN(\mult_49/ab[2][18] ), .OUT(n917) );
  INV U693 ( .IN(\mult_49/ab[3][17] ), .OUT(n918) );
  NAND2 U694 ( .A(n920), .B(n921), .OUT(n919) );
  INV U695 ( .IN(\mult_49/ab[4][16] ), .OUT(n922) );
  NAND2 U696 ( .A(n924), .B(n925), .OUT(n923) );
  INV U697 ( .IN(\mult_49/ab[5][15] ), .OUT(n926) );
  NAND2 U698 ( .A(n928), .B(n929), .OUT(n927) );
  INV U699 ( .IN(\mult_49/ab[6][14] ), .OUT(n930) );
  NAND2 U700 ( .A(n932), .B(n933), .OUT(n931) );
  INV U701 ( .IN(\mult_49/ab[7][13] ), .OUT(n934) );
  NAND2 U702 ( .A(n936), .B(n937), .OUT(n935) );
  INV U703 ( .IN(\mult_49/ab[8][12] ), .OUT(n938) );
  NAND2 U704 ( .A(n940), .B(n941), .OUT(n939) );
  INV U705 ( .IN(\mult_49/ab[9][11] ), .OUT(n942) );
  NAND2 U706 ( .A(n944), .B(n945), .OUT(n943) );
  INV U707 ( .IN(\mult_49/ab[10][10] ), .OUT(n946) );
  NAND2 U708 ( .A(n948), .B(n949), .OUT(n947) );
  INV U709 ( .IN(\mult_49/ab[11][9] ), .OUT(n950) );
  NAND2 U710 ( .A(n952), .B(n953), .OUT(n951) );
  INV U711 ( .IN(\mult_49/ab[12][8] ), .OUT(n954) );
  NAND2 U712 ( .A(n956), .B(n957), .OUT(n955) );
  INV U713 ( .IN(\mult_49/ab[13][7] ), .OUT(n958) );
  NAND2 U714 ( .A(n960), .B(n961), .OUT(n959) );
  INV U715 ( .IN(\mult_49/ab[14][6] ), .OUT(n962) );
  NAND2 U716 ( .A(n964), .B(n965), .OUT(n963) );
  INV U717 ( .IN(\mult_49/ab[15][5] ), .OUT(n966) );
  NAND2 U718 ( .A(n968), .B(n969), .OUT(n967) );
  INV U719 ( .IN(\mult_49/ab[16][4] ), .OUT(n970) );
  NAND2 U720 ( .A(n972), .B(n973), .OUT(n971) );
  INV U721 ( .IN(\mult_49/ab[17][3] ), .OUT(n974) );
  NAND2 U722 ( .A(n976), .B(n977), .OUT(n975) );
  INV U723 ( .IN(\mult_49/ab[18][2] ), .OUT(n978) );
  NAND2 U724 ( .A(n980), .B(n981), .OUT(n979) );
  NOR2 U725 ( .A(n983), .B(n984), .OUT(n982) );
  INV U726 ( .IN(\mult_49/ab[2][19] ), .OUT(n985) );
  INV U727 ( .IN(\mult_49/ab[3][18] ), .OUT(n986) );
  NAND2 U728 ( .A(n988), .B(n989), .OUT(n987) );
  INV U729 ( .IN(\mult_49/ab[4][17] ), .OUT(n990) );
  NAND2 U730 ( .A(n992), .B(n993), .OUT(n991) );
  INV U731 ( .IN(\mult_49/ab[5][16] ), .OUT(n994) );
  NAND2 U732 ( .A(n996), .B(n997), .OUT(n995) );
  INV U733 ( .IN(\mult_49/ab[6][15] ), .OUT(n998) );
  NAND2 U734 ( .A(n1000), .B(n1001), .OUT(n999) );
  INV U735 ( .IN(\mult_49/ab[7][14] ), .OUT(n1002) );
  NAND2 U736 ( .A(n1004), .B(n1005), .OUT(n1003) );
  INV U737 ( .IN(\mult_49/ab[8][13] ), .OUT(n1006) );
  NAND2 U738 ( .A(n1008), .B(n1009), .OUT(n1007) );
  INV U739 ( .IN(\mult_49/ab[9][12] ), .OUT(n1010) );
  NAND2 U740 ( .A(n1012), .B(n1013), .OUT(n1011) );
  INV U741 ( .IN(\mult_49/ab[10][11] ), .OUT(n1014) );
  NAND2 U742 ( .A(n1016), .B(n1017), .OUT(n1015) );
  INV U743 ( .IN(\mult_49/ab[11][10] ), .OUT(n1018) );
  NAND2 U744 ( .A(n1020), .B(n1021), .OUT(n1019) );
  INV U745 ( .IN(\mult_49/ab[12][9] ), .OUT(n1022) );
  NAND2 U746 ( .A(n1024), .B(n1025), .OUT(n1023) );
  INV U747 ( .IN(\mult_49/ab[13][8] ), .OUT(n1026) );
  NAND2 U748 ( .A(n1028), .B(n1029), .OUT(n1027) );
  INV U749 ( .IN(\mult_49/ab[14][7] ), .OUT(n1030) );
  NAND2 U750 ( .A(n1032), .B(n1033), .OUT(n1031) );
  INV U751 ( .IN(\mult_49/ab[15][6] ), .OUT(n1034) );
  NAND2 U752 ( .A(n1036), .B(n1037), .OUT(n1035) );
  INV U753 ( .IN(\mult_49/ab[16][5] ), .OUT(n1038) );
  NAND2 U754 ( .A(n1040), .B(n1041), .OUT(n1039) );
  INV U755 ( .IN(\mult_49/ab[17][4] ), .OUT(n1042) );
  NAND2 U756 ( .A(n1044), .B(n1045), .OUT(n1043) );
  INV U757 ( .IN(\mult_49/ab[18][3] ), .OUT(n1046) );
  NAND2 U758 ( .A(n1048), .B(n1049), .OUT(n1047) );
  INV U759 ( .IN(\mult_49/ab[19][2] ), .OUT(n1050) );
  NAND2 U760 ( .A(n1052), .B(n1053), .OUT(n1051) );
  NOR2 U761 ( .A(n1055), .B(n1056), .OUT(n1054) );
  INV U762 ( .IN(\mult_49/ab[2][20] ), .OUT(n1057) );
  INV U763 ( .IN(\mult_49/ab[3][19] ), .OUT(n1058) );
  NAND2 U764 ( .A(n1060), .B(n1061), .OUT(n1059) );
  INV U765 ( .IN(\mult_49/ab[4][18] ), .OUT(n1062) );
  NAND2 U766 ( .A(n1064), .B(n1065), .OUT(n1063) );
  INV U767 ( .IN(\mult_49/ab[5][17] ), .OUT(n1066) );
  NAND2 U768 ( .A(n1068), .B(n1069), .OUT(n1067) );
  INV U769 ( .IN(\mult_49/ab[6][16] ), .OUT(n1070) );
  NAND2 U770 ( .A(n1072), .B(n1073), .OUT(n1071) );
  INV U771 ( .IN(\mult_49/ab[7][15] ), .OUT(n1074) );
  NAND2 U772 ( .A(n1076), .B(n1077), .OUT(n1075) );
  INV U773 ( .IN(\mult_49/ab[8][14] ), .OUT(n1078) );
  NAND2 U774 ( .A(n1080), .B(n1081), .OUT(n1079) );
  INV U775 ( .IN(\mult_49/ab[9][13] ), .OUT(n1082) );
  NAND2 U776 ( .A(n1084), .B(n1085), .OUT(n1083) );
  INV U777 ( .IN(\mult_49/ab[10][12] ), .OUT(n1086) );
  NAND2 U778 ( .A(n1088), .B(n1089), .OUT(n1087) );
  INV U779 ( .IN(\mult_49/ab[11][11] ), .OUT(n1090) );
  NAND2 U780 ( .A(n1092), .B(n1093), .OUT(n1091) );
  INV U781 ( .IN(\mult_49/ab[12][10] ), .OUT(n1094) );
  NAND2 U782 ( .A(n1096), .B(n1097), .OUT(n1095) );
  INV U783 ( .IN(\mult_49/ab[13][9] ), .OUT(n1098) );
  NAND2 U784 ( .A(n1100), .B(n1101), .OUT(n1099) );
  INV U785 ( .IN(\mult_49/ab[14][8] ), .OUT(n1102) );
  NAND2 U786 ( .A(n1104), .B(n1105), .OUT(n1103) );
  INV U787 ( .IN(\mult_49/ab[15][7] ), .OUT(n1106) );
  NAND2 U788 ( .A(n1108), .B(n1109), .OUT(n1107) );
  INV U789 ( .IN(\mult_49/ab[16][6] ), .OUT(n1110) );
  NAND2 U790 ( .A(n1112), .B(n1113), .OUT(n1111) );
  INV U791 ( .IN(\mult_49/ab[17][5] ), .OUT(n1114) );
  NAND2 U792 ( .A(n1116), .B(n1117), .OUT(n1115) );
  INV U793 ( .IN(\mult_49/ab[18][4] ), .OUT(n1118) );
  NAND2 U794 ( .A(n1120), .B(n1121), .OUT(n1119) );
  INV U795 ( .IN(\mult_49/ab[19][3] ), .OUT(n1122) );
  NAND2 U796 ( .A(n1124), .B(n1125), .OUT(n1123) );
  INV U797 ( .IN(\mult_49/ab[20][2] ), .OUT(n1126) );
  NAND2 U798 ( .A(n1128), .B(n1129), .OUT(n1127) );
  NOR2 U799 ( .A(n1131), .B(n1132), .OUT(n1130) );
  INV U800 ( .IN(\mult_49/ab[2][21] ), .OUT(n1133) );
  INV U801 ( .IN(\mult_49/ab[3][20] ), .OUT(n1134) );
  NAND2 U802 ( .A(n1136), .B(n1137), .OUT(n1135) );
  INV U803 ( .IN(\mult_49/ab[4][19] ), .OUT(n1138) );
  NAND2 U804 ( .A(n1140), .B(n1141), .OUT(n1139) );
  INV U805 ( .IN(\mult_49/ab[5][18] ), .OUT(n1142) );
  NAND2 U806 ( .A(n1144), .B(n1145), .OUT(n1143) );
  INV U807 ( .IN(\mult_49/ab[6][17] ), .OUT(n1146) );
  NAND2 U808 ( .A(n1148), .B(n1149), .OUT(n1147) );
  INV U809 ( .IN(\mult_49/ab[7][16] ), .OUT(n1150) );
  NAND2 U810 ( .A(n1152), .B(n1153), .OUT(n1151) );
  INV U811 ( .IN(\mult_49/ab[8][15] ), .OUT(n1154) );
  NAND2 U812 ( .A(n1156), .B(n1157), .OUT(n1155) );
  INV U813 ( .IN(\mult_49/ab[9][14] ), .OUT(n1158) );
  NAND2 U814 ( .A(n1160), .B(n1161), .OUT(n1159) );
  INV U815 ( .IN(\mult_49/ab[10][13] ), .OUT(n1162) );
  NAND2 U816 ( .A(n1164), .B(n1165), .OUT(n1163) );
  INV U817 ( .IN(\mult_49/ab[11][12] ), .OUT(n1166) );
  NAND2 U818 ( .A(n1168), .B(n1169), .OUT(n1167) );
  INV U819 ( .IN(\mult_49/ab[12][11] ), .OUT(n1170) );
  NAND2 U820 ( .A(n1172), .B(n1173), .OUT(n1171) );
  INV U821 ( .IN(\mult_49/ab[13][10] ), .OUT(n1174) );
  NAND2 U822 ( .A(n1176), .B(n1177), .OUT(n1175) );
  INV U823 ( .IN(\mult_49/ab[14][9] ), .OUT(n1178) );
  NAND2 U824 ( .A(n1180), .B(n1181), .OUT(n1179) );
  INV U825 ( .IN(\mult_49/ab[15][8] ), .OUT(n1182) );
  NAND2 U826 ( .A(n1184), .B(n1185), .OUT(n1183) );
  INV U827 ( .IN(\mult_49/ab[16][7] ), .OUT(n1186) );
  NAND2 U828 ( .A(n1188), .B(n1189), .OUT(n1187) );
  INV U829 ( .IN(\mult_49/ab[17][6] ), .OUT(n1190) );
  NAND2 U830 ( .A(n1192), .B(n1193), .OUT(n1191) );
  INV U831 ( .IN(\mult_49/ab[18][5] ), .OUT(n1194) );
  NAND2 U832 ( .A(n1196), .B(n1197), .OUT(n1195) );
  INV U833 ( .IN(\mult_49/ab[19][4] ), .OUT(n1198) );
  NAND2 U834 ( .A(n1200), .B(n1201), .OUT(n1199) );
  INV U835 ( .IN(\mult_49/ab[20][3] ), .OUT(n1202) );
  NAND2 U836 ( .A(n1204), .B(n1205), .OUT(n1203) );
  INV U837 ( .IN(\mult_49/ab[21][2] ), .OUT(n1206) );
  NAND2 U838 ( .A(n1208), .B(n1209), .OUT(n1207) );
  NOR2 U839 ( .A(n1211), .B(n1212), .OUT(n1210) );
  INV U840 ( .IN(\mult_49/ab[2][22] ), .OUT(n1213) );
  INV U841 ( .IN(\mult_49/ab[3][21] ), .OUT(n1214) );
  NAND2 U842 ( .A(n1216), .B(n1217), .OUT(n1215) );
  INV U843 ( .IN(\mult_49/ab[4][20] ), .OUT(n1218) );
  NAND2 U844 ( .A(n1220), .B(n1221), .OUT(n1219) );
  INV U845 ( .IN(\mult_49/ab[5][19] ), .OUT(n1222) );
  NAND2 U846 ( .A(n1224), .B(n1225), .OUT(n1223) );
  INV U847 ( .IN(\mult_49/ab[6][18] ), .OUT(n1226) );
  NAND2 U848 ( .A(n1228), .B(n1229), .OUT(n1227) );
  INV U849 ( .IN(\mult_49/ab[7][17] ), .OUT(n1230) );
  NAND2 U850 ( .A(n1232), .B(n1233), .OUT(n1231) );
  INV U851 ( .IN(\mult_49/ab[8][16] ), .OUT(n1234) );
  NAND2 U852 ( .A(n1236), .B(n1237), .OUT(n1235) );
  INV U853 ( .IN(\mult_49/ab[9][15] ), .OUT(n1238) );
  NAND2 U854 ( .A(n1240), .B(n1241), .OUT(n1239) );
  INV U855 ( .IN(\mult_49/ab[10][14] ), .OUT(n1242) );
  NAND2 U856 ( .A(n1244), .B(n1245), .OUT(n1243) );
  INV U857 ( .IN(\mult_49/ab[11][13] ), .OUT(n1246) );
  NAND2 U858 ( .A(n1248), .B(n1249), .OUT(n1247) );
  INV U859 ( .IN(\mult_49/ab[12][12] ), .OUT(n1250) );
  NAND2 U860 ( .A(n1252), .B(n1253), .OUT(n1251) );
  INV U861 ( .IN(\mult_49/ab[13][11] ), .OUT(n1254) );
  NAND2 U862 ( .A(n1256), .B(n1257), .OUT(n1255) );
  INV U863 ( .IN(\mult_49/ab[14][10] ), .OUT(n1258) );
  NAND2 U864 ( .A(n1260), .B(n1261), .OUT(n1259) );
  INV U865 ( .IN(\mult_49/ab[15][9] ), .OUT(n1262) );
  NAND2 U866 ( .A(n1264), .B(n1265), .OUT(n1263) );
  INV U867 ( .IN(\mult_49/ab[16][8] ), .OUT(n1266) );
  NAND2 U868 ( .A(n1268), .B(n1269), .OUT(n1267) );
  INV U869 ( .IN(\mult_49/ab[17][7] ), .OUT(n1270) );
  NAND2 U870 ( .A(n1272), .B(n1273), .OUT(n1271) );
  INV U871 ( .IN(\mult_49/ab[18][6] ), .OUT(n1274) );
  NAND2 U872 ( .A(n1276), .B(n1277), .OUT(n1275) );
  INV U873 ( .IN(\mult_49/ab[19][5] ), .OUT(n1278) );
  NAND2 U874 ( .A(n1280), .B(n1281), .OUT(n1279) );
  INV U875 ( .IN(\mult_49/ab[20][4] ), .OUT(n1282) );
  NAND2 U876 ( .A(n1284), .B(n1285), .OUT(n1283) );
  INV U877 ( .IN(\mult_49/ab[21][3] ), .OUT(n1286) );
  NAND2 U878 ( .A(n1288), .B(n1289), .OUT(n1287) );
  INV U879 ( .IN(\mult_49/ab[22][2] ), .OUT(n1290) );
  NAND2 U880 ( .A(n1292), .B(n1293), .OUT(n1291) );
  NOR2 U881 ( .A(n1295), .B(n1296), .OUT(n1294) );
  INV U882 ( .IN(\mult_49/ab[2][23] ), .OUT(n1297) );
  INV U883 ( .IN(\mult_49/ab[3][22] ), .OUT(n1298) );
  NAND2 U884 ( .A(n1300), .B(n1301), .OUT(n1299) );
  INV U885 ( .IN(\mult_49/ab[4][21] ), .OUT(n1302) );
  NAND2 U886 ( .A(n1304), .B(n1305), .OUT(n1303) );
  INV U887 ( .IN(\mult_49/ab[5][20] ), .OUT(n1306) );
  NAND2 U888 ( .A(n1308), .B(n1309), .OUT(n1307) );
  INV U889 ( .IN(\mult_49/ab[6][19] ), .OUT(n1310) );
  NAND2 U890 ( .A(n1312), .B(n1313), .OUT(n1311) );
  INV U891 ( .IN(\mult_49/ab[7][18] ), .OUT(n1314) );
  NAND2 U892 ( .A(n1316), .B(n1317), .OUT(n1315) );
  INV U893 ( .IN(\mult_49/ab[8][17] ), .OUT(n1318) );
  NAND2 U894 ( .A(n1320), .B(n1321), .OUT(n1319) );
  INV U895 ( .IN(\mult_49/ab[9][16] ), .OUT(n1322) );
  NAND2 U896 ( .A(n1324), .B(n1325), .OUT(n1323) );
  INV U897 ( .IN(\mult_49/ab[10][15] ), .OUT(n1326) );
  NAND2 U898 ( .A(n1328), .B(n1329), .OUT(n1327) );
  INV U899 ( .IN(\mult_49/ab[11][14] ), .OUT(n1330) );
  NAND2 U900 ( .A(n1332), .B(n1333), .OUT(n1331) );
  INV U901 ( .IN(\mult_49/ab[12][13] ), .OUT(n1334) );
  NAND2 U902 ( .A(n1336), .B(n1337), .OUT(n1335) );
  INV U903 ( .IN(\mult_49/ab[13][12] ), .OUT(n1338) );
  NAND2 U904 ( .A(n1340), .B(n1341), .OUT(n1339) );
  INV U905 ( .IN(\mult_49/ab[14][11] ), .OUT(n1342) );
  NAND2 U906 ( .A(n1344), .B(n1345), .OUT(n1343) );
  INV U907 ( .IN(\mult_49/ab[15][10] ), .OUT(n1346) );
  NAND2 U908 ( .A(n1348), .B(n1349), .OUT(n1347) );
  INV U909 ( .IN(\mult_49/ab[16][9] ), .OUT(n1350) );
  NAND2 U910 ( .A(n1352), .B(n1353), .OUT(n1351) );
  INV U911 ( .IN(\mult_49/ab[17][8] ), .OUT(n1354) );
  NAND2 U912 ( .A(n1356), .B(n1357), .OUT(n1355) );
  INV U913 ( .IN(\mult_49/ab[18][7] ), .OUT(n1358) );
  NAND2 U914 ( .A(n1360), .B(n1361), .OUT(n1359) );
  INV U915 ( .IN(\mult_49/ab[19][6] ), .OUT(n1362) );
  NAND2 U916 ( .A(n1364), .B(n1365), .OUT(n1363) );
  INV U917 ( .IN(\mult_49/ab[20][5] ), .OUT(n1366) );
  NAND2 U918 ( .A(n1368), .B(n1369), .OUT(n1367) );
  INV U919 ( .IN(\mult_49/ab[21][4] ), .OUT(n1370) );
  NAND2 U920 ( .A(n1372), .B(n1373), .OUT(n1371) );
  INV U921 ( .IN(\mult_49/ab[22][3] ), .OUT(n1374) );
  NAND2 U922 ( .A(n1376), .B(n1377), .OUT(n1375) );
  INV U923 ( .IN(\mult_49/ab[23][2] ), .OUT(n1378) );
  NAND2 U924 ( .A(n1380), .B(n1381), .OUT(n1379) );
  NOR2 U925 ( .A(n1383), .B(n1384), .OUT(n1382) );
  INV U926 ( .IN(\mult_49/ab[2][24] ), .OUT(n1385) );
  INV U927 ( .IN(\mult_49/ab[3][23] ), .OUT(n1386) );
  NAND2 U928 ( .A(n1388), .B(n1389), .OUT(n1387) );
  INV U929 ( .IN(\mult_49/ab[4][22] ), .OUT(n1390) );
  NAND2 U930 ( .A(n1392), .B(n1393), .OUT(n1391) );
  INV U931 ( .IN(\mult_49/ab[5][21] ), .OUT(n1394) );
  NAND2 U932 ( .A(n1396), .B(n1397), .OUT(n1395) );
  INV U933 ( .IN(\mult_49/ab[6][20] ), .OUT(n1398) );
  NAND2 U934 ( .A(n1400), .B(n1401), .OUT(n1399) );
  INV U935 ( .IN(\mult_49/ab[7][19] ), .OUT(n1402) );
  NAND2 U936 ( .A(n1404), .B(n1405), .OUT(n1403) );
  INV U937 ( .IN(\mult_49/ab[8][18] ), .OUT(n1406) );
  NAND2 U938 ( .A(n1408), .B(n1409), .OUT(n1407) );
  INV U939 ( .IN(\mult_49/ab[9][17] ), .OUT(n1410) );
  NAND2 U940 ( .A(n1412), .B(n1413), .OUT(n1411) );
  INV U941 ( .IN(\mult_49/ab[10][16] ), .OUT(n1414) );
  NAND2 U942 ( .A(n1416), .B(n1417), .OUT(n1415) );
  INV U943 ( .IN(\mult_49/ab[11][15] ), .OUT(n1418) );
  NAND2 U944 ( .A(n1420), .B(n1421), .OUT(n1419) );
  INV U945 ( .IN(\mult_49/ab[12][14] ), .OUT(n1422) );
  NAND2 U946 ( .A(n1424), .B(n1425), .OUT(n1423) );
  INV U947 ( .IN(\mult_49/ab[13][13] ), .OUT(n1426) );
  NAND2 U948 ( .A(n1428), .B(n1429), .OUT(n1427) );
  INV U949 ( .IN(\mult_49/ab[14][12] ), .OUT(n1430) );
  NAND2 U950 ( .A(n1432), .B(n1433), .OUT(n1431) );
  INV U951 ( .IN(\mult_49/ab[15][11] ), .OUT(n1434) );
  NAND2 U952 ( .A(n1436), .B(n1437), .OUT(n1435) );
  INV U953 ( .IN(\mult_49/ab[16][10] ), .OUT(n1438) );
  NAND2 U954 ( .A(n1440), .B(n1441), .OUT(n1439) );
  INV U955 ( .IN(\mult_49/ab[17][9] ), .OUT(n1442) );
  NAND2 U956 ( .A(n1444), .B(n1445), .OUT(n1443) );
  INV U957 ( .IN(\mult_49/ab[18][8] ), .OUT(n1446) );
  NAND2 U958 ( .A(n1448), .B(n1449), .OUT(n1447) );
  INV U959 ( .IN(\mult_49/ab[19][7] ), .OUT(n1450) );
  NAND2 U960 ( .A(n1452), .B(n1453), .OUT(n1451) );
  INV U961 ( .IN(\mult_49/ab[20][6] ), .OUT(n1454) );
  NAND2 U962 ( .A(n1456), .B(n1457), .OUT(n1455) );
  INV U963 ( .IN(\mult_49/ab[21][5] ), .OUT(n1458) );
  NAND2 U964 ( .A(n1460), .B(n1461), .OUT(n1459) );
  INV U965 ( .IN(\mult_49/ab[22][4] ), .OUT(n1462) );
  NAND2 U966 ( .A(n1464), .B(n1465), .OUT(n1463) );
  INV U967 ( .IN(\mult_49/ab[23][3] ), .OUT(n1466) );
  NAND2 U968 ( .A(n1468), .B(n1469), .OUT(n1467) );
  INV U969 ( .IN(\mult_49/ab[24][2] ), .OUT(n1470) );
  NAND2 U970 ( .A(n1472), .B(n1473), .OUT(n1471) );
  NOR2 U971 ( .A(n1475), .B(n1476), .OUT(n1474) );
  INV U972 ( .IN(\mult_49/ab[2][25] ), .OUT(n1477) );
  INV U973 ( .IN(\mult_49/ab[3][24] ), .OUT(n1478) );
  NAND2 U974 ( .A(n1480), .B(n1481), .OUT(n1479) );
  INV U975 ( .IN(\mult_49/ab[4][23] ), .OUT(n1482) );
  NAND2 U976 ( .A(n1484), .B(n1485), .OUT(n1483) );
  INV U977 ( .IN(\mult_49/ab[5][22] ), .OUT(n1486) );
  NAND2 U978 ( .A(n1488), .B(n1489), .OUT(n1487) );
  INV U979 ( .IN(\mult_49/ab[6][21] ), .OUT(n1490) );
  NAND2 U980 ( .A(n1492), .B(n1493), .OUT(n1491) );
  INV U981 ( .IN(\mult_49/ab[7][20] ), .OUT(n1494) );
  NAND2 U982 ( .A(n1496), .B(n1497), .OUT(n1495) );
  INV U983 ( .IN(\mult_49/ab[8][19] ), .OUT(n1498) );
  NAND2 U984 ( .A(n1500), .B(n1501), .OUT(n1499) );
  INV U985 ( .IN(\mult_49/ab[9][18] ), .OUT(n1502) );
  NAND2 U986 ( .A(n1504), .B(n1505), .OUT(n1503) );
  INV U987 ( .IN(\mult_49/ab[10][17] ), .OUT(n1506) );
  NAND2 U988 ( .A(n1508), .B(n1509), .OUT(n1507) );
  INV U989 ( .IN(\mult_49/ab[11][16] ), .OUT(n1510) );
  NAND2 U990 ( .A(n1512), .B(n1513), .OUT(n1511) );
  INV U991 ( .IN(\mult_49/ab[12][15] ), .OUT(n1514) );
  NAND2 U992 ( .A(n1516), .B(n1517), .OUT(n1515) );
  INV U993 ( .IN(\mult_49/ab[13][14] ), .OUT(n1518) );
  NAND2 U994 ( .A(n1520), .B(n1521), .OUT(n1519) );
  INV U995 ( .IN(\mult_49/ab[14][13] ), .OUT(n1522) );
  NAND2 U996 ( .A(n1524), .B(n1525), .OUT(n1523) );
  INV U997 ( .IN(\mult_49/ab[15][12] ), .OUT(n1526) );
  NAND2 U998 ( .A(n1528), .B(n1529), .OUT(n1527) );
  INV U999 ( .IN(\mult_49/ab[16][11] ), .OUT(n1530) );
  NAND2 U1000 ( .A(n1532), .B(n1533), .OUT(n1531) );
  INV U1001 ( .IN(\mult_49/ab[17][10] ), .OUT(n1534) );
  NAND2 U1002 ( .A(n1536), .B(n1537), .OUT(n1535) );
  INV U1003 ( .IN(\mult_49/ab[18][9] ), .OUT(n1538) );
  NAND2 U1004 ( .A(n1540), .B(n1541), .OUT(n1539) );
  INV U1005 ( .IN(\mult_49/ab[19][8] ), .OUT(n1542) );
  NAND2 U1006 ( .A(n1544), .B(n1545), .OUT(n1543) );
  INV U1007 ( .IN(\mult_49/ab[20][7] ), .OUT(n1546) );
  NAND2 U1008 ( .A(n1548), .B(n1549), .OUT(n1547) );
  INV U1009 ( .IN(\mult_49/ab[21][6] ), .OUT(n1550) );
  NAND2 U1010 ( .A(n1552), .B(n1553), .OUT(n1551) );
  INV U1011 ( .IN(\mult_49/ab[22][5] ), .OUT(n1554) );
  NAND2 U1012 ( .A(n1556), .B(n1557), .OUT(n1555) );
  INV U1013 ( .IN(\mult_49/ab[23][4] ), .OUT(n1558) );
  NAND2 U1014 ( .A(n1560), .B(n1561), .OUT(n1559) );
  INV U1015 ( .IN(\mult_49/ab[24][3] ), .OUT(n1562) );
  NAND2 U1016 ( .A(n1564), .B(n1565), .OUT(n1563) );
  INV U1017 ( .IN(\mult_49/ab[25][2] ), .OUT(n1566) );
  NAND2 U1018 ( .A(n1568), .B(n1569), .OUT(n1567) );
  NOR2 U1019 ( .A(n1571), .B(n1572), .OUT(n1570) );
  INV U1020 ( .IN(\mult_49/ab[2][26] ), .OUT(n1573) );
  INV U1021 ( .IN(\mult_49/ab[3][25] ), .OUT(n1574) );
  NAND2 U1022 ( .A(n1576), .B(n1577), .OUT(n1575) );
  INV U1023 ( .IN(\mult_49/ab[4][24] ), .OUT(n1578) );
  NAND2 U1024 ( .A(n1580), .B(n1581), .OUT(n1579) );
  INV U1025 ( .IN(\mult_49/ab[5][23] ), .OUT(n1582) );
  NAND2 U1026 ( .A(n1584), .B(n1585), .OUT(n1583) );
  INV U1027 ( .IN(\mult_49/ab[6][22] ), .OUT(n1586) );
  NAND2 U1028 ( .A(n1588), .B(n1589), .OUT(n1587) );
  INV U1029 ( .IN(\mult_49/ab[7][21] ), .OUT(n1590) );
  NAND2 U1030 ( .A(n1592), .B(n1593), .OUT(n1591) );
  INV U1031 ( .IN(\mult_49/ab[8][20] ), .OUT(n1594) );
  NAND2 U1032 ( .A(n1596), .B(n1597), .OUT(n1595) );
  INV U1033 ( .IN(\mult_49/ab[9][19] ), .OUT(n1598) );
  NAND2 U1034 ( .A(n1600), .B(n1601), .OUT(n1599) );
  INV U1035 ( .IN(\mult_49/ab[10][18] ), .OUT(n1602) );
  NAND2 U1036 ( .A(n1604), .B(n1605), .OUT(n1603) );
  INV U1037 ( .IN(\mult_49/ab[11][17] ), .OUT(n1606) );
  NAND2 U1038 ( .A(n1608), .B(n1609), .OUT(n1607) );
  INV U1039 ( .IN(\mult_49/ab[12][16] ), .OUT(n1610) );
  NAND2 U1040 ( .A(n1612), .B(n1613), .OUT(n1611) );
  INV U1041 ( .IN(\mult_49/ab[13][15] ), .OUT(n1614) );
  NAND2 U1042 ( .A(n1616), .B(n1617), .OUT(n1615) );
  INV U1043 ( .IN(\mult_49/ab[14][14] ), .OUT(n1618) );
  NAND2 U1044 ( .A(n1620), .B(n1621), .OUT(n1619) );
  INV U1045 ( .IN(\mult_49/ab[15][13] ), .OUT(n1622) );
  NAND2 U1046 ( .A(n1624), .B(n1625), .OUT(n1623) );
  INV U1047 ( .IN(\mult_49/ab[16][12] ), .OUT(n1626) );
  NAND2 U1048 ( .A(n1628), .B(n1629), .OUT(n1627) );
  INV U1049 ( .IN(\mult_49/ab[17][11] ), .OUT(n1630) );
  NAND2 U1050 ( .A(n1632), .B(n1633), .OUT(n1631) );
  INV U1051 ( .IN(\mult_49/ab[18][10] ), .OUT(n1634) );
  NAND2 U1052 ( .A(n1636), .B(n1637), .OUT(n1635) );
  INV U1053 ( .IN(\mult_49/ab[19][9] ), .OUT(n1638) );
  NAND2 U1054 ( .A(n1640), .B(n1641), .OUT(n1639) );
  INV U1055 ( .IN(\mult_49/ab[20][8] ), .OUT(n1642) );
  NAND2 U1056 ( .A(n1644), .B(n1645), .OUT(n1643) );
  INV U1057 ( .IN(\mult_49/ab[21][7] ), .OUT(n1646) );
  NAND2 U1058 ( .A(n1648), .B(n1649), .OUT(n1647) );
  INV U1059 ( .IN(\mult_49/ab[22][6] ), .OUT(n1650) );
  NAND2 U1060 ( .A(n1652), .B(n1653), .OUT(n1651) );
  INV U1061 ( .IN(\mult_49/ab[23][5] ), .OUT(n1654) );
  NAND2 U1062 ( .A(n1656), .B(n1657), .OUT(n1655) );
  INV U1063 ( .IN(\mult_49/ab[24][4] ), .OUT(n1658) );
  NAND2 U1064 ( .A(n1660), .B(n1661), .OUT(n1659) );
  INV U1065 ( .IN(\mult_49/ab[25][3] ), .OUT(n1662) );
  NAND2 U1066 ( .A(n1664), .B(n1665), .OUT(n1663) );
  INV U1067 ( .IN(\mult_49/ab[26][2] ), .OUT(n1666) );
  NAND2 U1068 ( .A(n1668), .B(n1669), .OUT(n1667) );
  NOR2 U1069 ( .A(n1671), .B(n1672), .OUT(n1670) );
  INV U1070 ( .IN(\mult_49/ab[2][27] ), .OUT(n1673) );
  INV U1071 ( .IN(\mult_49/ab[3][26] ), .OUT(n1674) );
  NAND2 U1072 ( .A(n1676), .B(n1677), .OUT(n1675) );
  INV U1073 ( .IN(\mult_49/ab[4][25] ), .OUT(n1678) );
  NAND2 U1074 ( .A(n1680), .B(n1681), .OUT(n1679) );
  INV U1075 ( .IN(\mult_49/ab[5][24] ), .OUT(n1682) );
  NAND2 U1076 ( .A(n1684), .B(n1685), .OUT(n1683) );
  INV U1077 ( .IN(\mult_49/ab[6][23] ), .OUT(n1686) );
  NAND2 U1078 ( .A(n1688), .B(n1689), .OUT(n1687) );
  INV U1079 ( .IN(\mult_49/ab[7][22] ), .OUT(n1690) );
  NAND2 U1080 ( .A(n1692), .B(n1693), .OUT(n1691) );
  INV U1081 ( .IN(\mult_49/ab[8][21] ), .OUT(n1694) );
  NAND2 U1082 ( .A(n1696), .B(n1697), .OUT(n1695) );
  INV U1083 ( .IN(\mult_49/ab[9][20] ), .OUT(n1698) );
  NAND2 U1084 ( .A(n1700), .B(n1701), .OUT(n1699) );
  INV U1085 ( .IN(\mult_49/ab[10][19] ), .OUT(n1702) );
  NAND2 U1086 ( .A(n1704), .B(n1705), .OUT(n1703) );
  INV U1087 ( .IN(\mult_49/ab[11][18] ), .OUT(n1706) );
  NAND2 U1088 ( .A(n1708), .B(n1709), .OUT(n1707) );
  INV U1089 ( .IN(\mult_49/ab[12][17] ), .OUT(n1710) );
  NAND2 U1090 ( .A(n1712), .B(n1713), .OUT(n1711) );
  INV U1091 ( .IN(\mult_49/ab[13][16] ), .OUT(n1714) );
  NAND2 U1092 ( .A(n1716), .B(n1717), .OUT(n1715) );
  INV U1093 ( .IN(\mult_49/ab[14][15] ), .OUT(n1718) );
  NAND2 U1094 ( .A(n1720), .B(n1721), .OUT(n1719) );
  INV U1095 ( .IN(\mult_49/ab[15][14] ), .OUT(n1722) );
  NAND2 U1096 ( .A(n1724), .B(n1725), .OUT(n1723) );
  INV U1097 ( .IN(\mult_49/ab[16][13] ), .OUT(n1726) );
  NAND2 U1098 ( .A(n1728), .B(n1729), .OUT(n1727) );
  INV U1099 ( .IN(\mult_49/ab[17][12] ), .OUT(n1730) );
  NAND2 U1100 ( .A(n1732), .B(n1733), .OUT(n1731) );
  INV U1101 ( .IN(\mult_49/ab[18][11] ), .OUT(n1734) );
  NAND2 U1102 ( .A(n1736), .B(n1737), .OUT(n1735) );
  INV U1103 ( .IN(\mult_49/ab[19][10] ), .OUT(n1738) );
  NAND2 U1104 ( .A(n1740), .B(n1741), .OUT(n1739) );
  INV U1105 ( .IN(\mult_49/ab[20][9] ), .OUT(n1742) );
  NAND2 U1106 ( .A(n1744), .B(n1745), .OUT(n1743) );
  INV U1107 ( .IN(\mult_49/ab[21][8] ), .OUT(n1746) );
  NAND2 U1108 ( .A(n1748), .B(n1749), .OUT(n1747) );
  INV U1109 ( .IN(\mult_49/ab[22][7] ), .OUT(n1750) );
  NAND2 U1110 ( .A(n1752), .B(n1753), .OUT(n1751) );
  INV U1111 ( .IN(\mult_49/ab[23][6] ), .OUT(n1754) );
  NAND2 U1112 ( .A(n1756), .B(n1757), .OUT(n1755) );
  INV U1113 ( .IN(\mult_49/ab[24][5] ), .OUT(n1758) );
  NAND2 U1114 ( .A(n1760), .B(n1761), .OUT(n1759) );
  INV U1115 ( .IN(\mult_49/ab[25][4] ), .OUT(n1762) );
  NAND2 U1116 ( .A(n1764), .B(n1765), .OUT(n1763) );
  INV U1117 ( .IN(\mult_49/ab[26][3] ), .OUT(n1766) );
  NAND2 U1118 ( .A(n1768), .B(n1769), .OUT(n1767) );
  INV U1119 ( .IN(\mult_49/ab[27][2] ), .OUT(n1770) );
  NAND2 U1120 ( .A(n1772), .B(n1773), .OUT(n1771) );
  NOR2 U1121 ( .A(n1775), .B(n1776), .OUT(n1774) );
  INV U1122 ( .IN(\mult_49/ab[2][28] ), .OUT(n1777) );
  INV U1123 ( .IN(\mult_49/ab[3][27] ), .OUT(n1778) );
  NAND2 U1124 ( .A(n1780), .B(n1781), .OUT(n1779) );
  INV U1125 ( .IN(\mult_49/ab[4][26] ), .OUT(n1782) );
  NAND2 U1126 ( .A(n1784), .B(n1785), .OUT(n1783) );
  INV U1127 ( .IN(\mult_49/ab[5][25] ), .OUT(n1786) );
  NAND2 U1128 ( .A(n1788), .B(n1789), .OUT(n1787) );
  INV U1129 ( .IN(\mult_49/ab[6][24] ), .OUT(n1790) );
  NAND2 U1130 ( .A(n1792), .B(n1793), .OUT(n1791) );
  INV U1131 ( .IN(\mult_49/ab[7][23] ), .OUT(n1794) );
  NAND2 U1132 ( .A(n1796), .B(n1797), .OUT(n1795) );
  INV U1133 ( .IN(\mult_49/ab[8][22] ), .OUT(n1798) );
  NAND2 U1134 ( .A(n1800), .B(n1801), .OUT(n1799) );
  INV U1135 ( .IN(\mult_49/ab[9][21] ), .OUT(n1802) );
  NAND2 U1136 ( .A(n1804), .B(n1805), .OUT(n1803) );
  INV U1137 ( .IN(\mult_49/ab[10][20] ), .OUT(n1806) );
  NAND2 U1138 ( .A(n1808), .B(n1809), .OUT(n1807) );
  INV U1139 ( .IN(\mult_49/ab[11][19] ), .OUT(n1810) );
  NAND2 U1140 ( .A(n1812), .B(n1813), .OUT(n1811) );
  INV U1141 ( .IN(\mult_49/ab[12][18] ), .OUT(n1814) );
  NAND2 U1142 ( .A(n1816), .B(n1817), .OUT(n1815) );
  INV U1143 ( .IN(\mult_49/ab[13][17] ), .OUT(n1818) );
  NAND2 U1144 ( .A(n1820), .B(n1821), .OUT(n1819) );
  INV U1145 ( .IN(\mult_49/ab[14][16] ), .OUT(n1822) );
  NAND2 U1146 ( .A(n1824), .B(n1825), .OUT(n1823) );
  INV U1147 ( .IN(\mult_49/ab[15][15] ), .OUT(n1826) );
  NAND2 U1148 ( .A(n1828), .B(n1829), .OUT(n1827) );
  INV U1149 ( .IN(\mult_49/ab[16][14] ), .OUT(n1830) );
  NAND2 U1150 ( .A(n1832), .B(n1833), .OUT(n1831) );
  INV U1151 ( .IN(\mult_49/ab[17][13] ), .OUT(n1834) );
  NAND2 U1152 ( .A(n1836), .B(n1837), .OUT(n1835) );
  INV U1153 ( .IN(\mult_49/ab[18][12] ), .OUT(n1838) );
  NAND2 U1154 ( .A(n1840), .B(n1841), .OUT(n1839) );
  INV U1155 ( .IN(\mult_49/ab[19][11] ), .OUT(n1842) );
  NAND2 U1156 ( .A(n1844), .B(n1845), .OUT(n1843) );
  INV U1157 ( .IN(\mult_49/ab[20][10] ), .OUT(n1846) );
  NAND2 U1158 ( .A(n1848), .B(n1849), .OUT(n1847) );
  INV U1159 ( .IN(\mult_49/ab[21][9] ), .OUT(n1850) );
  NAND2 U1160 ( .A(n1852), .B(n1853), .OUT(n1851) );
  INV U1161 ( .IN(\mult_49/ab[22][8] ), .OUT(n1854) );
  NAND2 U1162 ( .A(n1856), .B(n1857), .OUT(n1855) );
  INV U1163 ( .IN(\mult_49/ab[23][7] ), .OUT(n1858) );
  NAND2 U1164 ( .A(n1860), .B(n1861), .OUT(n1859) );
  INV U1165 ( .IN(\mult_49/ab[24][6] ), .OUT(n1862) );
  NAND2 U1166 ( .A(n1864), .B(n1865), .OUT(n1863) );
  INV U1167 ( .IN(\mult_49/ab[25][5] ), .OUT(n1866) );
  NAND2 U1168 ( .A(n1868), .B(n1869), .OUT(n1867) );
  INV U1169 ( .IN(\mult_49/ab[26][4] ), .OUT(n1870) );
  NAND2 U1170 ( .A(n1872), .B(n1873), .OUT(n1871) );
  INV U1171 ( .IN(\mult_49/ab[27][3] ), .OUT(n1874) );
  NAND2 U1172 ( .A(n1876), .B(n1877), .OUT(n1875) );
  INV U1173 ( .IN(\mult_49/ab[28][2] ), .OUT(n1878) );
  NAND2 U1174 ( .A(n1880), .B(n1881), .OUT(n1879) );
  INV U1175 ( .IN(\mult_49/ab[11][1] ), .OUT(n1882) );
  NAND2 U1176 ( .A(n1884), .B(n1885), .OUT(n1883) );
  INV U1177 ( .IN(\mult_49/ab[12][1] ), .OUT(n1886) );
  NAND2 U1178 ( .A(n1888), .B(n1889), .OUT(n1887) );
  INV U1179 ( .IN(\mult_49/ab[13][1] ), .OUT(n1890) );
  NAND2 U1180 ( .A(n1892), .B(n1893), .OUT(n1891) );
  INV U1181 ( .IN(\mult_49/ab[14][1] ), .OUT(n1894) );
  NAND2 U1182 ( .A(n1896), .B(n1897), .OUT(n1895) );
  INV U1183 ( .IN(\mult_49/ab[15][1] ), .OUT(n1898) );
  NAND2 U1184 ( .A(n1900), .B(n1901), .OUT(n1899) );
  INV U1185 ( .IN(\mult_49/ab[16][1] ), .OUT(n1902) );
  NAND2 U1186 ( .A(n1904), .B(n1905), .OUT(n1903) );
  INV U1187 ( .IN(\mult_49/ab[17][1] ), .OUT(n1906) );
  NAND2 U1188 ( .A(n1908), .B(n1909), .OUT(n1907) );
  INV U1189 ( .IN(\mult_49/ab[18][1] ), .OUT(n1910) );
  NAND2 U1190 ( .A(n1912), .B(n1913), .OUT(n1911) );
  INV U1191 ( .IN(\mult_49/ab[19][1] ), .OUT(n1914) );
  NAND2 U1192 ( .A(n1916), .B(n1917), .OUT(n1915) );
  INV U1193 ( .IN(\mult_49/ab[20][1] ), .OUT(n1918) );
  NAND2 U1194 ( .A(n1920), .B(n1921), .OUT(n1919) );
  INV U1195 ( .IN(\mult_49/ab[21][1] ), .OUT(n1922) );
  NAND2 U1196 ( .A(n1924), .B(n1925), .OUT(n1923) );
  INV U1197 ( .IN(\mult_49/ab[22][1] ), .OUT(n1926) );
  NAND2 U1198 ( .A(n1928), .B(n1929), .OUT(n1927) );
  INV U1199 ( .IN(\mult_49/ab[23][1] ), .OUT(n1930) );
  NAND2 U1200 ( .A(n1932), .B(n1933), .OUT(n1931) );
  INV U1201 ( .IN(\mult_49/ab[24][1] ), .OUT(n1934) );
  NAND2 U1202 ( .A(n1936), .B(n1937), .OUT(n1935) );
  INV U1203 ( .IN(\mult_49/ab[25][1] ), .OUT(n1938) );
  NAND2 U1204 ( .A(n1940), .B(n1941), .OUT(n1939) );
  INV U1205 ( .IN(\mult_49/ab[26][1] ), .OUT(n1942) );
  NAND2 U1206 ( .A(n1944), .B(n1945), .OUT(n1943) );
  INV U1207 ( .IN(\mult_49/ab[27][1] ), .OUT(n1946) );
  NAND2 U1208 ( .A(n1948), .B(n1949), .OUT(n1947) );
  INV U1209 ( .IN(\mult_49/ab[28][1] ), .OUT(n1950) );
  NAND2 U1210 ( .A(n1952), .B(n1953), .OUT(n1951) );
  INV U1211 ( .IN(\mult_49/ab[29][1] ), .OUT(n1954) );
  NAND2 U1212 ( .A(n1956), .B(n1957), .OUT(n1955) );
  INV U1213 ( .IN(\mult_49/ab[12][0] ), .OUT(n1958) );
  NAND2 U1214 ( .A(n1960), .B(n1961), .OUT(n1959) );
  INV U1215 ( .IN(\mult_49/ab[13][0] ), .OUT(n1962) );
  NAND2 U1216 ( .A(n1964), .B(n1965), .OUT(n1963) );
  INV U1217 ( .IN(\mult_49/ab[14][0] ), .OUT(n1966) );
  NAND2 U1218 ( .A(n1968), .B(n1969), .OUT(n1967) );
  INV U1219 ( .IN(\mult_49/ab[15][0] ), .OUT(n1970) );
  NAND2 U1220 ( .A(n1972), .B(n1973), .OUT(n1971) );
  INV U1221 ( .IN(\mult_49/ab[16][0] ), .OUT(n1974) );
  NAND2 U1222 ( .A(n1976), .B(n1977), .OUT(n1975) );
  INV U1223 ( .IN(\mult_49/ab[17][0] ), .OUT(n1978) );
  NAND2 U1224 ( .A(n1980), .B(n1981), .OUT(n1979) );
  INV U1225 ( .IN(\mult_49/ab[18][0] ), .OUT(n1982) );
  NAND2 U1226 ( .A(n1984), .B(n1985), .OUT(n1983) );
  INV U1227 ( .IN(\mult_49/ab[19][0] ), .OUT(n1986) );
  NAND2 U1228 ( .A(n1988), .B(n1989), .OUT(n1987) );
  INV U1229 ( .IN(\mult_49/ab[20][0] ), .OUT(n1990) );
  NAND2 U1230 ( .A(n1992), .B(n1993), .OUT(n1991) );
  INV U1231 ( .IN(\mult_49/ab[21][0] ), .OUT(n1994) );
  NAND2 U1232 ( .A(n1996), .B(n1997), .OUT(n1995) );
  INV U1233 ( .IN(\mult_49/ab[22][0] ), .OUT(n1998) );
  NAND2 U1234 ( .A(n2000), .B(n2001), .OUT(n1999) );
  INV U1235 ( .IN(\mult_49/ab[23][0] ), .OUT(n2002) );
  NAND2 U1236 ( .A(n2004), .B(n2005), .OUT(n2003) );
  INV U1237 ( .IN(\mult_49/ab[24][0] ), .OUT(n2006) );
  NAND2 U1238 ( .A(n2008), .B(n2009), .OUT(n2007) );
  INV U1239 ( .IN(\mult_49/ab[25][0] ), .OUT(n2010) );
  NAND2 U1240 ( .A(n2012), .B(n2013), .OUT(n2011) );
  INV U1241 ( .IN(\mult_49/ab[26][0] ), .OUT(n2014) );
  NAND2 U1242 ( .A(n2016), .B(n2017), .OUT(n2015) );
  INV U1243 ( .IN(\mult_49/ab[27][0] ), .OUT(n2018) );
  NAND2 U1244 ( .A(n2020), .B(n2021), .OUT(n2019) );
  INV U1245 ( .IN(\mult_49/ab[28][0] ), .OUT(n2022) );
  NAND2 U1246 ( .A(n2024), .B(n2025), .OUT(n2023) );
  INV U1247 ( .IN(\mult_49/ab[29][0] ), .OUT(n2026) );
  NAND2 U1248 ( .A(n2028), .B(n2029), .OUT(n2027) );
  INV U1249 ( .IN(\mult_49/ab[30][0] ), .OUT(n2030) );
  INV U1250 ( .IN(A[9]), .OUT(n2031) );
  INV U1251 ( .IN(B[9]), .OUT(n2032) );
  INV U1252 ( .IN(A[8]), .OUT(n2033) );
  INV U1253 ( .IN(B[8]), .OUT(n2034) );
  INV U1254 ( .IN(A[7]), .OUT(n2035) );
  INV U1255 ( .IN(B[7]), .OUT(n2036) );
  INV U1256 ( .IN(A[6]), .OUT(n2037) );
  INV U1257 ( .IN(B[6]), .OUT(n2038) );
  INV U1258 ( .IN(A[5]), .OUT(n2039) );
  INV U1259 ( .IN(B[5]), .OUT(n2040) );
  INV U1260 ( .IN(A[4]), .OUT(n2041) );
  INV U1261 ( .IN(B[4]), .OUT(n2042) );
  INV U1262 ( .IN(A[3]), .OUT(n2043) );
  INV U1263 ( .IN(B[3]), .OUT(n2044) );
  INV U1264 ( .IN(A[30]), .OUT(n2045) );
  INV U1265 ( .IN(B[30]), .OUT(n2046) );
  INV U1266 ( .IN(A[2]), .OUT(n2047) );
  INV U1267 ( .IN(B[2]), .OUT(n2048) );
  INV U1268 ( .IN(A[29]), .OUT(n2049) );
  INV U1269 ( .IN(B[29]), .OUT(n2050) );
  INV U1270 ( .IN(A[28]), .OUT(n2051) );
  INV U1271 ( .IN(B[28]), .OUT(n2052) );
  INV U1272 ( .IN(A[27]), .OUT(n2053) );
  INV U1273 ( .IN(B[27]), .OUT(n2054) );
  INV U1274 ( .IN(A[26]), .OUT(n2055) );
  INV U1275 ( .IN(B[26]), .OUT(n2056) );
  INV U1276 ( .IN(A[25]), .OUT(n2057) );
  INV U1277 ( .IN(B[25]), .OUT(n2058) );
  INV U1278 ( .IN(A[24]), .OUT(n2059) );
  INV U1279 ( .IN(B[24]), .OUT(n2060) );
  INV U1280 ( .IN(A[23]), .OUT(n2061) );
  INV U1281 ( .IN(B[23]), .OUT(n2062) );
  INV U1282 ( .IN(A[22]), .OUT(n2063) );
  INV U1283 ( .IN(B[22]), .OUT(n2064) );
  INV U1284 ( .IN(A[21]), .OUT(n2065) );
  INV U1285 ( .IN(B[21]), .OUT(n2066) );
  INV U1286 ( .IN(A[20]), .OUT(n2067) );
  INV U1287 ( .IN(B[20]), .OUT(n2068) );
  INV U1288 ( .IN(A[1]), .OUT(n2069) );
  INV U1289 ( .IN(B[1]), .OUT(n2070) );
  INV U1290 ( .IN(A[19]), .OUT(n2071) );
  INV U1291 ( .IN(B[19]), .OUT(n2072) );
  INV U1292 ( .IN(A[18]), .OUT(n2073) );
  INV U1293 ( .IN(B[18]), .OUT(n2074) );
  INV U1294 ( .IN(A[17]), .OUT(n2075) );
  INV U1295 ( .IN(B[17]), .OUT(n2076) );
  INV U1296 ( .IN(A[16]), .OUT(n2077) );
  INV U1297 ( .IN(B[16]), .OUT(n2078) );
  INV U1298 ( .IN(A[15]), .OUT(n2079) );
  INV U1299 ( .IN(B[15]), .OUT(n2080) );
  INV U1300 ( .IN(A[14]), .OUT(n2081) );
  INV U1301 ( .IN(B[14]), .OUT(n2082) );
  INV U1302 ( .IN(A[13]), .OUT(n2083) );
  INV U1303 ( .IN(B[13]), .OUT(n2084) );
  INV U1304 ( .IN(A[12]), .OUT(n2085) );
  INV U1305 ( .IN(B[12]), .OUT(n2086) );
  INV U1306 ( .IN(A[11]), .OUT(n2087) );
  INV U1307 ( .IN(B[11]), .OUT(n2088) );
  INV U1308 ( .IN(A[10]), .OUT(n2089) );
  INV U1309 ( .IN(B[10]), .OUT(n2090) );
  NOR2 U1310 ( .A(\mult_49/A_notx[0] ), .B(\mult_49/B_notx[0] ), .OUT(n2091)
         );
  NOR2 U1311 ( .A(\mult_49/B_notx[0] ), .B(A[0]), .OUT(n2092) );
  NAND2 U1312 ( .A(n2094), .B(n2095), .OUT(n2093) );
  NAND2 U1313 ( .A(n2097), .B(n2098), .OUT(n2096) );
  NAND2 U1314 ( .A(n2100), .B(n2101), .OUT(n2099) );
  NAND2 U1315 ( .A(n2103), .B(n2104), .OUT(n2102) );
  NAND2 U1316 ( .A(n2106), .B(n2107), .OUT(n2105) );
  NAND2 U1317 ( .A(n2109), .B(n2110), .OUT(n2108) );
  NAND2 U1318 ( .A(n2112), .B(n2113), .OUT(n2111) );
  NAND2 U1319 ( .A(n2115), .B(n2116), .OUT(n2114) );
  NAND2 U1320 ( .A(n2118), .B(n2119), .OUT(n2117) );
  NAND2 U1321 ( .A(n2121), .B(n2122), .OUT(n2120) );
  NAND2 U1322 ( .A(n2124), .B(n2125), .OUT(n2123) );
  NAND2 U1323 ( .A(n2127), .B(n2128), .OUT(n2126) );
  NAND2 U1324 ( .A(n2130), .B(n2131), .OUT(n2129) );
  NAND2 U1325 ( .A(n2133), .B(n2134), .OUT(n2132) );
  NAND2 U1326 ( .A(n2136), .B(n2137), .OUT(n2135) );
  NAND2 U1327 ( .A(n2139), .B(n2140), .OUT(n2138) );
  NAND2 U1328 ( .A(n2142), .B(n2143), .OUT(n2141) );
  NAND2 U1329 ( .A(n2145), .B(n2146), .OUT(n2144) );
  NAND2 U1330 ( .A(n2148), .B(n2149), .OUT(n2147) );
  NAND2 U1331 ( .A(n2151), .B(n2152), .OUT(n2150) );
  NAND2 U1332 ( .A(n2154), .B(n2155), .OUT(n2153) );
  NAND2 U1333 ( .A(n2157), .B(n2158), .OUT(n2156) );
  NAND2 U1334 ( .A(n2160), .B(n2161), .OUT(n2159) );
  NAND2 U1335 ( .A(n2163), .B(n2164), .OUT(n2162) );
  NAND2 U1336 ( .A(n2166), .B(n2167), .OUT(n2165) );
  NAND2 U1337 ( .A(n2169), .B(n2170), .OUT(n2168) );
  NAND2 U1338 ( .A(n2172), .B(n2173), .OUT(n2171) );
  NAND2 U1339 ( .A(n2175), .B(n2176), .OUT(n2174) );
  NAND2 U1340 ( .A(n2178), .B(n2179), .OUT(n2177) );
  NAND2 U1341 ( .A(n2181), .B(n2182), .OUT(n2180) );
  NAND2 U1342 ( .A(n2184), .B(n2185), .OUT(n2183) );
  NAND2 U1343 ( .A(n2187), .B(n2188), .OUT(n2186) );
  NOR2 U1344 ( .A(n2190), .B(n2191), .OUT(n2189) );
  NAND2 U1345 ( .A(n2193), .B(n2194), .OUT(n2192) );
  NAND2 U1346 ( .A(n2196), .B(n2197), .OUT(n2195) );
  NAND2 U1347 ( .A(n2199), .B(n2200), .OUT(n2198) );
  NAND2 U1348 ( .A(n2202), .B(n2203), .OUT(n2201) );
  NAND2 U1349 ( .A(n2205), .B(n2206), .OUT(n2204) );
  NOR2 U1350 ( .A(n2208), .B(n2209), .OUT(n2207) );
  NOR2 U1351 ( .A(n2211), .B(n2212), .OUT(n2210) );
  NAND2 U1352 ( .A(n2214), .B(n2215), .OUT(n2213) );
  NAND2 U1353 ( .A(n2217), .B(n2218), .OUT(n2216) );
  NOR2 U1354 ( .A(n2220), .B(n2221), .OUT(n2219) );
  NAND2 U1355 ( .A(n2223), .B(n2224), .OUT(n2222) );
  NAND2 U1356 ( .A(n2226), .B(n2227), .OUT(n2225) );
  NAND2 U1357 ( .A(n2229), .B(n2230), .OUT(n2228) );
  NAND2 U1358 ( .A(n2232), .B(n2233), .OUT(n2231) );
  NOR2 U1359 ( .A(n2235), .B(n2236), .OUT(n2234) );
  NAND2 U1360 ( .A(n2238), .B(n2239), .OUT(n2237) );
  NOR2 U1361 ( .A(n2241), .B(n2242), .OUT(n2240) );
  NOR2 U1362 ( .A(n2244), .B(n2245), .OUT(n2243) );
  NAND2 U1363 ( .A(n2247), .B(n2248), .OUT(n2246) );
  NAND2 U1364 ( .A(n2250), .B(n2251), .OUT(n2249) );
  NOR2 U1365 ( .A(n2253), .B(n2254), .OUT(n2252) );
  NAND2 U1366 ( .A(n2256), .B(n2257), .OUT(n2255) );
  NOR2 U1367 ( .A(n2259), .B(n2260), .OUT(n2258) );
  NAND2 U1368 ( .A(n2262), .B(n2263), .OUT(n2261) );
  NAND2 U1369 ( .A(n2265), .B(n2266), .OUT(n2264) );
  NAND2 U1370 ( .A(n2268), .B(n2269), .OUT(n2267) );
  NAND2 U1371 ( .A(n2271), .B(n2272), .OUT(n2270) );
  NOR2 U1372 ( .A(n2274), .B(n2275), .OUT(n2273) );
  NAND2 U1373 ( .A(n2277), .B(n2278), .OUT(n2276) );
  NOR2 U1374 ( .A(n2280), .B(n2281), .OUT(n2279) );
  NAND2 U1375 ( .A(n2283), .B(n2284), .OUT(n2282) );
  NOR2 U1376 ( .A(n2286), .B(n2287), .OUT(n2285) );
  NOR2 U1377 ( .A(n2289), .B(n2290), .OUT(n2288) );
  NAND2 U1378 ( .A(n2292), .B(n2293), .OUT(n2291) );
  NAND2 U1379 ( .A(n2295), .B(n2296), .OUT(n2294) );
  NOR2 U1380 ( .A(n2298), .B(n2299), .OUT(n2297) );
  NAND2 U1381 ( .A(n2301), .B(n2302), .OUT(n2300) );
  NOR2 U1382 ( .A(n2304), .B(n2305), .OUT(n2303) );
  NAND2 U1383 ( .A(n2307), .B(n2308), .OUT(n2306) );
  NOR2 U1384 ( .A(n2310), .B(n2311), .OUT(n2309) );
  NAND2 U1385 ( .A(n2313), .B(n2314), .OUT(n2312) );
  NOR2 U1386 ( .A(n2316), .B(n2317), .OUT(n2315) );
  NAND2 U1387 ( .A(n2319), .B(n2320), .OUT(n2318) );
  NOR2 U1388 ( .A(n2322), .B(n2323), .OUT(n2321) );
  NOR2 U1389 ( .A(n2325), .B(n2326), .OUT(n2324) );
  NOR2 U1390 ( .A(n2328), .B(n2329), .OUT(n2327) );
  NOR2 U1391 ( .A(n2331), .B(n2332), .OUT(n2330) );
  NOR2 U1392 ( .A(n2334), .B(n2335), .OUT(n2333) );
  NOR2 U1393 ( .A(n2337), .B(n2338), .OUT(n2336) );
  NOR2 U1394 ( .A(n2340), .B(n2341), .OUT(n2339) );
  NOR2 U1395 ( .A(n2343), .B(n2344), .OUT(n2342) );
  NAND2 U1396 ( .A(n2345), .B(n2346), .OUT(\mult_49/A1[8] ) );
  NAND2 U1397 ( .A(n2347), .B(n2348), .OUT(\mult_49/A1[6] ) );
  NAND2 U1398 ( .A(n2349), .B(n2350), .OUT(\mult_49/A1[4] ) );
  NAND2 U1399 ( .A(n2351), .B(n2352), .OUT(\mult_49/A1[2] ) );
  NAND2 U1400 ( .A(n2354), .B(n2355), .OUT(n2353) );
  NAND2 U1401 ( .A(n2357), .B(n2358), .OUT(n2356) );
  NOR2 U1402 ( .A(n2360), .B(n2361), .OUT(n2359) );
  NAND2 U1403 ( .A(n2363), .B(n2364), .OUT(n2362) );
  NOR2 U1404 ( .A(n2366), .B(n2367), .OUT(n2365) );
  NAND2 U1405 ( .A(n2369), .B(n2370), .OUT(n2368) );
  NOR2 U1406 ( .A(n2372), .B(n2373), .OUT(n2371) );
  NAND2 U1407 ( .A(n2375), .B(n2376), .OUT(n2374) );
  NOR2 U1408 ( .A(n2378), .B(n2379), .OUT(n2377) );
  NAND2 U1409 ( .A(n2381), .B(n2382), .OUT(n2380) );
  NAND2 U1410 ( .A(n2384), .B(n2385), .OUT(n2383) );
  NOR2 U1411 ( .A(n2387), .B(n2388), .OUT(n2386) );
  NAND2 U1412 ( .A(n2390), .B(n2391), .OUT(n2389) );
  NOR2 U1413 ( .A(n2393), .B(n2394), .OUT(n2392) );
  NAND2 U1414 ( .A(n2396), .B(n2397), .OUT(n2395) );
  NOR2 U1415 ( .A(n2399), .B(n2400), .OUT(n2398) );
  NAND2 U1416 ( .A(n2402), .B(n2403), .OUT(n2401) );
  NOR2 U1417 ( .A(n2405), .B(n2406), .OUT(n2404) );
  NAND2 U1418 ( .A(n2408), .B(n2409), .OUT(n2407) );
  NAND2 U1419 ( .A(n2411), .B(n2412), .OUT(n2410) );
  NAND2 U1420 ( .A(n2414), .B(n2415), .OUT(n2413) );
  NOR2 U1421 ( .A(n2417), .B(n2418), .OUT(n2416) );
  NAND2 U1422 ( .A(n2420), .B(n2421), .OUT(n2419) );
  NOR2 U1423 ( .A(n2423), .B(n2424), .OUT(n2422) );
  NAND2 U1424 ( .A(n2426), .B(n2427), .OUT(n2425) );
  NOR2 U1425 ( .A(n2429), .B(n2430), .OUT(n2428) );
  NAND2 U1426 ( .A(n2432), .B(n2433), .OUT(n2431) );
  NOR2 U1427 ( .A(n2435), .B(n2436), .OUT(n2434) );
  NAND2 U1428 ( .A(n2438), .B(n2439), .OUT(n2437) );
  NOR2 U1429 ( .A(n2441), .B(n2442), .OUT(n2440) );
  NAND2 U1430 ( .A(n2444), .B(n2445), .OUT(n2443) );
  NAND2 U1431 ( .A(n2447), .B(n2448), .OUT(n2446) );
  NOR2 U1432 ( .A(n2450), .B(n2451), .OUT(n2449) );
  NAND2 U1433 ( .A(n2453), .B(n2454), .OUT(n2452) );
  NOR2 U1434 ( .A(n2456), .B(n2457), .OUT(n2455) );
  NAND2 U1435 ( .A(n2459), .B(n2460), .OUT(n2458) );
  NOR2 U1436 ( .A(n2462), .B(n2463), .OUT(n2461) );
  NAND2 U1437 ( .A(n2465), .B(n2466), .OUT(n2464) );
  NOR2 U1438 ( .A(n2468), .B(n2469), .OUT(n2467) );
  NAND2 U1439 ( .A(n2471), .B(n2472), .OUT(n2470) );
  NOR2 U1440 ( .A(n2474), .B(n2475), .OUT(n2473) );
  NAND2 U1441 ( .A(n2477), .B(n2478), .OUT(n2476) );
  NAND2 U1442 ( .A(n2480), .B(n2481), .OUT(n2479) );
  NAND2 U1443 ( .A(n2483), .B(n2484), .OUT(n2482) );
  NOR2 U1444 ( .A(n2486), .B(n2487), .OUT(n2485) );
  NAND2 U1445 ( .A(n2489), .B(n2490), .OUT(n2488) );
  NOR2 U1446 ( .A(n2492), .B(n2493), .OUT(n2491) );
  NAND2 U1447 ( .A(n2495), .B(n2496), .OUT(n2494) );
  NOR2 U1448 ( .A(n2498), .B(n2499), .OUT(n2497) );
  NAND2 U1449 ( .A(n2501), .B(n2502), .OUT(n2500) );
  NOR2 U1450 ( .A(n2504), .B(n2505), .OUT(n2503) );
  NAND2 U1451 ( .A(n2507), .B(n2508), .OUT(n2506) );
  NOR2 U1452 ( .A(n2510), .B(n2511), .OUT(n2509) );
  NAND2 U1453 ( .A(n2513), .B(n2514), .OUT(n2512) );
  NOR2 U1454 ( .A(n2516), .B(n2517), .OUT(n2515) );
  NAND2 U1455 ( .A(n2519), .B(n2520), .OUT(n2518) );
  NAND2 U1456 ( .A(n2522), .B(n2523), .OUT(n2521) );
  NOR2 U1457 ( .A(n2525), .B(n2526), .OUT(n2524) );
  NAND2 U1458 ( .A(n2528), .B(n2529), .OUT(n2527) );
  NOR2 U1459 ( .A(n2531), .B(n2532), .OUT(n2530) );
  NAND2 U1460 ( .A(n2534), .B(n2535), .OUT(n2533) );
  NOR2 U1461 ( .A(n2537), .B(n2538), .OUT(n2536) );
  NAND2 U1462 ( .A(n2540), .B(n2541), .OUT(n2539) );
  NOR2 U1463 ( .A(n2543), .B(n2544), .OUT(n2542) );
  NAND2 U1464 ( .A(n2546), .B(n2547), .OUT(n2545) );
  NOR2 U1465 ( .A(n2549), .B(n2550), .OUT(n2548) );
  NAND2 U1466 ( .A(n2552), .B(n2553), .OUT(n2551) );
  NOR2 U1467 ( .A(n2555), .B(n2556), .OUT(n2554) );
  NAND2 U1468 ( .A(n2558), .B(n2559), .OUT(n2557) );
  NAND2 U1469 ( .A(n2561), .B(n2562), .OUT(n2560) );
  NAND2 U1470 ( .A(n2564), .B(n2565), .OUT(n2563) );
  NOR2 U1471 ( .A(n2567), .B(n2568), .OUT(n2566) );
  NAND2 U1472 ( .A(n2570), .B(n2571), .OUT(n2569) );
  NOR2 U1473 ( .A(n2573), .B(n2574), .OUT(n2572) );
  NAND2 U1474 ( .A(n2576), .B(n2577), .OUT(n2575) );
  NOR2 U1475 ( .A(n2579), .B(n2580), .OUT(n2578) );
  NAND2 U1476 ( .A(n2582), .B(n2583), .OUT(n2581) );
  NOR2 U1477 ( .A(n2585), .B(n2586), .OUT(n2584) );
  NAND2 U1478 ( .A(n2588), .B(n2589), .OUT(n2587) );
  NOR2 U1479 ( .A(n2591), .B(n2592), .OUT(n2590) );
  NAND2 U1480 ( .A(n2594), .B(n2595), .OUT(n2593) );
  NOR2 U1481 ( .A(n2597), .B(n2598), .OUT(n2596) );
  NAND2 U1482 ( .A(n2600), .B(n2601), .OUT(n2599) );
  NOR2 U1483 ( .A(n2603), .B(n2604), .OUT(n2602) );
  NAND2 U1484 ( .A(n2606), .B(n2607), .OUT(n2605) );
  NAND2 U1485 ( .A(n2609), .B(n2610), .OUT(n2608) );
  NOR2 U1486 ( .A(n2612), .B(n2613), .OUT(n2611) );
  NAND2 U1487 ( .A(n2615), .B(n2616), .OUT(n2614) );
  NOR2 U1488 ( .A(n2618), .B(n2619), .OUT(n2617) );
  NAND2 U1489 ( .A(n2621), .B(n2622), .OUT(n2620) );
  NOR2 U1490 ( .A(n2624), .B(n2625), .OUT(n2623) );
  NAND2 U1491 ( .A(n2627), .B(n2628), .OUT(n2626) );
  NOR2 U1492 ( .A(n2630), .B(n2631), .OUT(n2629) );
  NAND2 U1493 ( .A(n2633), .B(n2634), .OUT(n2632) );
  NOR2 U1494 ( .A(n2636), .B(n2637), .OUT(n2635) );
  NAND2 U1495 ( .A(n2639), .B(n2640), .OUT(n2638) );
  NOR2 U1496 ( .A(n2642), .B(n2643), .OUT(n2641) );
  NAND2 U1497 ( .A(n2645), .B(n2646), .OUT(n2644) );
  NOR2 U1498 ( .A(n2648), .B(n2649), .OUT(n2647) );
  NAND2 U1499 ( .A(n2651), .B(n2652), .OUT(n2650) );
  NAND2 U1500 ( .A(n2654), .B(n2655), .OUT(n2653) );
  NAND2 U1501 ( .A(n2657), .B(n2658), .OUT(n2656) );
  NOR2 U1502 ( .A(n2660), .B(n2661), .OUT(n2659) );
  NAND2 U1503 ( .A(n2663), .B(n2664), .OUT(n2662) );
  NOR2 U1504 ( .A(n2666), .B(n2667), .OUT(n2665) );
  NAND2 U1505 ( .A(n2669), .B(n2670), .OUT(n2668) );
  NOR2 U1506 ( .A(n2672), .B(n2673), .OUT(n2671) );
  NAND2 U1507 ( .A(n2675), .B(n2676), .OUT(n2674) );
  NOR2 U1508 ( .A(n2678), .B(n2679), .OUT(n2677) );
  NAND2 U1509 ( .A(n2681), .B(n2682), .OUT(n2680) );
  NOR2 U1510 ( .A(n2684), .B(n2685), .OUT(n2683) );
  NAND2 U1511 ( .A(n2687), .B(n2688), .OUT(n2686) );
  NOR2 U1512 ( .A(n2690), .B(n2691), .OUT(n2689) );
  NAND2 U1513 ( .A(n2693), .B(n2694), .OUT(n2692) );
  NOR2 U1514 ( .A(n2696), .B(n2697), .OUT(n2695) );
  NAND2 U1515 ( .A(n2699), .B(n2700), .OUT(n2698) );
  NOR2 U1516 ( .A(n2702), .B(n2703), .OUT(n2701) );
  NAND2 U1517 ( .A(n2705), .B(n2706), .OUT(n2704) );
  NAND2 U1518 ( .A(n2708), .B(n2709), .OUT(n2707) );
  NOR2 U1519 ( .A(n2711), .B(n2712), .OUT(n2710) );
  NAND2 U1520 ( .A(n2714), .B(n2715), .OUT(n2713) );
  NOR2 U1521 ( .A(n2717), .B(n2718), .OUT(n2716) );
  NAND2 U1522 ( .A(n2720), .B(n2721), .OUT(n2719) );
  NOR2 U1523 ( .A(n2723), .B(n2724), .OUT(n2722) );
  NAND2 U1524 ( .A(n2726), .B(n2727), .OUT(n2725) );
  NOR2 U1525 ( .A(n2729), .B(n2730), .OUT(n2728) );
  NAND2 U1526 ( .A(n2732), .B(n2733), .OUT(n2731) );
  NOR2 U1527 ( .A(n2735), .B(n2736), .OUT(n2734) );
  NAND2 U1528 ( .A(n2738), .B(n2739), .OUT(n2737) );
  NOR2 U1529 ( .A(n2741), .B(n2742), .OUT(n2740) );
  NAND2 U1530 ( .A(n2744), .B(n2745), .OUT(n2743) );
  NOR2 U1531 ( .A(n2747), .B(n2748), .OUT(n2746) );
  NAND2 U1532 ( .A(n2750), .B(n2751), .OUT(n2749) );
  NOR2 U1533 ( .A(n2753), .B(n2754), .OUT(n2752) );
  NAND2 U1534 ( .A(n2756), .B(n2757), .OUT(n2755) );
  NAND2 U1535 ( .A(n2759), .B(n2760), .OUT(n2758) );
  NAND2 U1536 ( .A(n2762), .B(n2763), .OUT(n2761) );
  NOR2 U1537 ( .A(n2765), .B(n2766), .OUT(n2764) );
  NAND2 U1538 ( .A(n2768), .B(n2769), .OUT(n2767) );
  NOR2 U1539 ( .A(n2771), .B(n2772), .OUT(n2770) );
  NAND2 U1540 ( .A(n2774), .B(n2775), .OUT(n2773) );
  NOR2 U1541 ( .A(n2777), .B(n2778), .OUT(n2776) );
  NAND2 U1542 ( .A(n2780), .B(n2781), .OUT(n2779) );
  NOR2 U1543 ( .A(n2783), .B(n2784), .OUT(n2782) );
  NAND2 U1544 ( .A(n2786), .B(n2787), .OUT(n2785) );
  NOR2 U1545 ( .A(n2789), .B(n2790), .OUT(n2788) );
  NAND2 U1546 ( .A(n2792), .B(n2793), .OUT(n2791) );
  NOR2 U1547 ( .A(n2795), .B(n2796), .OUT(n2794) );
  NAND2 U1548 ( .A(n2798), .B(n2799), .OUT(n2797) );
  NOR2 U1549 ( .A(n2801), .B(n2802), .OUT(n2800) );
  NAND2 U1550 ( .A(n2804), .B(n2805), .OUT(n2803) );
  NOR2 U1551 ( .A(n2807), .B(n2808), .OUT(n2806) );
  NAND2 U1552 ( .A(n2810), .B(n2811), .OUT(n2809) );
  NOR2 U1553 ( .A(n2813), .B(n2814), .OUT(n2812) );
  NAND2 U1554 ( .A(n2816), .B(n2817), .OUT(n2815) );
  NAND2 U1555 ( .A(n2819), .B(n2820), .OUT(n2818) );
  NOR2 U1556 ( .A(n2822), .B(n2823), .OUT(n2821) );
  NAND2 U1557 ( .A(n2825), .B(n2826), .OUT(n2824) );
  NOR2 U1558 ( .A(n2828), .B(n2829), .OUT(n2827) );
  NAND2 U1559 ( .A(n2831), .B(n2832), .OUT(n2830) );
  NOR2 U1560 ( .A(n2834), .B(n2835), .OUT(n2833) );
  NAND2 U1561 ( .A(n2837), .B(n2838), .OUT(n2836) );
  NOR2 U1562 ( .A(n2840), .B(n2841), .OUT(n2839) );
  NAND2 U1563 ( .A(n2843), .B(n2844), .OUT(n2842) );
  NOR2 U1564 ( .A(n2846), .B(n2847), .OUT(n2845) );
  NAND2 U1565 ( .A(n2849), .B(n2850), .OUT(n2848) );
  NOR2 U1566 ( .A(n2852), .B(n2853), .OUT(n2851) );
  NAND2 U1567 ( .A(n2855), .B(n2856), .OUT(n2854) );
  NOR2 U1568 ( .A(n2858), .B(n2859), .OUT(n2857) );
  NAND2 U1569 ( .A(n2861), .B(n2862), .OUT(n2860) );
  NOR2 U1570 ( .A(n2864), .B(n2865), .OUT(n2863) );
  NAND2 U1571 ( .A(n2867), .B(n2868), .OUT(n2866) );
  NOR2 U1572 ( .A(n2870), .B(n2871), .OUT(n2869) );
  NAND2 U1573 ( .A(n2873), .B(n2874), .OUT(n2872) );
  NAND2 U1574 ( .A(n2876), .B(n2877), .OUT(n2875) );
  NAND2 U1575 ( .A(n2879), .B(n2880), .OUT(n2878) );
  NOR2 U1576 ( .A(n2882), .B(n2883), .OUT(n2881) );
  NAND2 U1577 ( .A(n2885), .B(n2886), .OUT(n2884) );
  NOR2 U1578 ( .A(n2888), .B(n2889), .OUT(n2887) );
  NAND2 U1579 ( .A(n2891), .B(n2892), .OUT(n2890) );
  NOR2 U1580 ( .A(n2894), .B(n2895), .OUT(n2893) );
  NAND2 U1581 ( .A(n2897), .B(n2898), .OUT(n2896) );
  NOR2 U1582 ( .A(n2900), .B(n2901), .OUT(n2899) );
  NAND2 U1583 ( .A(n2903), .B(n2904), .OUT(n2902) );
  NOR2 U1584 ( .A(n2906), .B(n2907), .OUT(n2905) );
  NAND2 U1585 ( .A(n2909), .B(n2910), .OUT(n2908) );
  NOR2 U1586 ( .A(n2912), .B(n2913), .OUT(n2911) );
  NAND2 U1587 ( .A(n2915), .B(n2916), .OUT(n2914) );
  NOR2 U1588 ( .A(n2918), .B(n2919), .OUT(n2917) );
  NAND2 U1589 ( .A(n2921), .B(n2922), .OUT(n2920) );
  NOR2 U1590 ( .A(n2924), .B(n2925), .OUT(n2923) );
  NAND2 U1591 ( .A(n2927), .B(n2928), .OUT(n2926) );
  NOR2 U1592 ( .A(n2930), .B(n2931), .OUT(n2929) );
  NAND2 U1593 ( .A(n2933), .B(n2934), .OUT(n2932) );
  NOR2 U1594 ( .A(n2936), .B(n2937), .OUT(n2935) );
  NAND2 U1595 ( .A(n2939), .B(n2940), .OUT(n2938) );
  NAND2 U1596 ( .A(n2942), .B(n2943), .OUT(n2941) );
  NOR2 U1597 ( .A(n2945), .B(n2946), .OUT(n2944) );
  NAND2 U1598 ( .A(n2948), .B(n2949), .OUT(n2947) );
  NOR2 U1599 ( .A(n2951), .B(n2952), .OUT(n2950) );
  NAND2 U1600 ( .A(n2954), .B(n2955), .OUT(n2953) );
  NOR2 U1601 ( .A(n2957), .B(n2958), .OUT(n2956) );
  NAND2 U1602 ( .A(n2960), .B(n2961), .OUT(n2959) );
  NOR2 U1603 ( .A(n2963), .B(n2964), .OUT(n2962) );
  NAND2 U1604 ( .A(n2966), .B(n2967), .OUT(n2965) );
  NOR2 U1605 ( .A(n2969), .B(n2970), .OUT(n2968) );
  NAND2 U1606 ( .A(n2972), .B(n2973), .OUT(n2971) );
  NOR2 U1607 ( .A(n2975), .B(n2976), .OUT(n2974) );
  NAND2 U1608 ( .A(n2978), .B(n2979), .OUT(n2977) );
  NOR2 U1609 ( .A(n2981), .B(n2982), .OUT(n2980) );
  NAND2 U1610 ( .A(n2984), .B(n2985), .OUT(n2983) );
  NOR2 U1611 ( .A(n2987), .B(n2988), .OUT(n2986) );
  NAND2 U1612 ( .A(n2990), .B(n2991), .OUT(n2989) );
  NOR2 U1613 ( .A(n2993), .B(n2994), .OUT(n2992) );
  NAND2 U1614 ( .A(n2996), .B(n2997), .OUT(n2995) );
  NOR2 U1615 ( .A(n2999), .B(n3000), .OUT(n2998) );
  NAND2 U1616 ( .A(n3002), .B(n3003), .OUT(n3001) );
  NAND2 U1617 ( .A(n3005), .B(n3006), .OUT(n3004) );
  NAND2 U1618 ( .A(n3008), .B(n3009), .OUT(n3007) );
  NOR2 U1619 ( .A(n3011), .B(n3012), .OUT(n3010) );
  NAND2 U1620 ( .A(n3014), .B(n3015), .OUT(n3013) );
  NOR2 U1621 ( .A(n3017), .B(n3018), .OUT(n3016) );
  NAND2 U1622 ( .A(n3020), .B(n3021), .OUT(n3019) );
  NOR2 U1623 ( .A(n3023), .B(n3024), .OUT(n3022) );
  NAND2 U1624 ( .A(n3026), .B(n3027), .OUT(n3025) );
  NOR2 U1625 ( .A(n3029), .B(n3030), .OUT(n3028) );
  NAND2 U1626 ( .A(n3032), .B(n3033), .OUT(n3031) );
  NOR2 U1627 ( .A(n3035), .B(n3036), .OUT(n3034) );
  NAND2 U1628 ( .A(n3038), .B(n3039), .OUT(n3037) );
  NOR2 U1629 ( .A(n3041), .B(n3042), .OUT(n3040) );
  NAND2 U1630 ( .A(n3044), .B(n3045), .OUT(n3043) );
  NOR2 U1631 ( .A(n3047), .B(n3048), .OUT(n3046) );
  NAND2 U1632 ( .A(n3050), .B(n3051), .OUT(n3049) );
  NOR2 U1633 ( .A(n3053), .B(n3054), .OUT(n3052) );
  NAND2 U1634 ( .A(n3056), .B(n3057), .OUT(n3055) );
  NOR2 U1635 ( .A(n3059), .B(n3060), .OUT(n3058) );
  NAND2 U1636 ( .A(n3062), .B(n3063), .OUT(n3061) );
  NOR2 U1637 ( .A(n3065), .B(n3066), .OUT(n3064) );
  NAND2 U1638 ( .A(n3068), .B(n3069), .OUT(n3067) );
  NOR2 U1639 ( .A(n3071), .B(n3072), .OUT(n3070) );
  NAND2 U1640 ( .A(n3074), .B(n3075), .OUT(n3073) );
  NAND2 U1641 ( .A(n3077), .B(n3078), .OUT(n3076) );
  NOR2 U1642 ( .A(n3080), .B(n3081), .OUT(n3079) );
  NAND2 U1643 ( .A(n3083), .B(n3084), .OUT(n3082) );
  NOR2 U1644 ( .A(n3086), .B(n3087), .OUT(n3085) );
  NAND2 U1645 ( .A(n3089), .B(n3090), .OUT(n3088) );
  NOR2 U1646 ( .A(n3092), .B(n3093), .OUT(n3091) );
  NAND2 U1647 ( .A(n3095), .B(n3096), .OUT(n3094) );
  NOR2 U1648 ( .A(n3098), .B(n3099), .OUT(n3097) );
  NAND2 U1649 ( .A(n3101), .B(n3102), .OUT(n3100) );
  NOR2 U1650 ( .A(n3104), .B(n3105), .OUT(n3103) );
  NAND2 U1651 ( .A(n3107), .B(n3108), .OUT(n3106) );
  NOR2 U1652 ( .A(n3110), .B(n3111), .OUT(n3109) );
  NAND2 U1653 ( .A(n3113), .B(n3114), .OUT(n3112) );
  NOR2 U1654 ( .A(n3116), .B(n3117), .OUT(n3115) );
  NAND2 U1655 ( .A(n3119), .B(n3120), .OUT(n3118) );
  NOR2 U1656 ( .A(n3122), .B(n3123), .OUT(n3121) );
  NAND2 U1657 ( .A(n3125), .B(n3126), .OUT(n3124) );
  NOR2 U1658 ( .A(n3128), .B(n3129), .OUT(n3127) );
  NAND2 U1659 ( .A(n3131), .B(n3132), .OUT(n3130) );
  NOR2 U1660 ( .A(n3134), .B(n3135), .OUT(n3133) );
  NAND2 U1661 ( .A(n3137), .B(n3138), .OUT(n3136) );
  NOR2 U1662 ( .A(n3140), .B(n3141), .OUT(n3139) );
  NAND2 U1663 ( .A(n3143), .B(n3144), .OUT(n3142) );
  NAND2 U1664 ( .A(n3146), .B(n3147), .OUT(n3145) );
  NAND2 U1665 ( .A(n3149), .B(n3150), .OUT(n3148) );
  NOR2 U1666 ( .A(n3152), .B(n3153), .OUT(n3151) );
  NAND2 U1667 ( .A(n3155), .B(n3156), .OUT(n3154) );
  NOR2 U1668 ( .A(n3158), .B(n3159), .OUT(n3157) );
  NAND2 U1669 ( .A(n3161), .B(n3162), .OUT(n3160) );
  NOR2 U1670 ( .A(n3164), .B(n3165), .OUT(n3163) );
  NAND2 U1671 ( .A(n3167), .B(n3168), .OUT(n3166) );
  NOR2 U1672 ( .A(n3170), .B(n3171), .OUT(n3169) );
  NAND2 U1673 ( .A(n3173), .B(n3174), .OUT(n3172) );
  NOR2 U1674 ( .A(n3176), .B(n3177), .OUT(n3175) );
  NAND2 U1675 ( .A(n3179), .B(n3180), .OUT(n3178) );
  NOR2 U1676 ( .A(n3182), .B(n3183), .OUT(n3181) );
  NAND2 U1677 ( .A(n3185), .B(n3186), .OUT(n3184) );
  NOR2 U1678 ( .A(n3188), .B(n3189), .OUT(n3187) );
  NAND2 U1679 ( .A(n3191), .B(n3192), .OUT(n3190) );
  NOR2 U1680 ( .A(n3194), .B(n3195), .OUT(n3193) );
  NAND2 U1681 ( .A(n3197), .B(n3198), .OUT(n3196) );
  NOR2 U1682 ( .A(n3200), .B(n3201), .OUT(n3199) );
  NAND2 U1683 ( .A(n3203), .B(n3204), .OUT(n3202) );
  NOR2 U1684 ( .A(n3206), .B(n3207), .OUT(n3205) );
  NAND2 U1685 ( .A(n3209), .B(n3210), .OUT(n3208) );
  NOR2 U1686 ( .A(n3212), .B(n3213), .OUT(n3211) );
  NAND2 U1687 ( .A(n3215), .B(n3216), .OUT(n3214) );
  NOR2 U1688 ( .A(n3218), .B(n3219), .OUT(n3217) );
  NAND2 U1689 ( .A(n3221), .B(n3222), .OUT(n3220) );
  NAND2 U1690 ( .A(n3224), .B(n3225), .OUT(n3223) );
  NOR2 U1691 ( .A(n3227), .B(n3228), .OUT(n3226) );
  NAND2 U1692 ( .A(n3230), .B(n3231), .OUT(n3229) );
  NOR2 U1693 ( .A(n3233), .B(n3234), .OUT(n3232) );
  NAND2 U1694 ( .A(n3236), .B(n3237), .OUT(n3235) );
  NOR2 U1695 ( .A(n3239), .B(n3240), .OUT(n3238) );
  NAND2 U1696 ( .A(n3242), .B(n3243), .OUT(n3241) );
  NOR2 U1697 ( .A(n3245), .B(n3246), .OUT(n3244) );
  NAND2 U1698 ( .A(n3248), .B(n3249), .OUT(n3247) );
  NOR2 U1699 ( .A(n3251), .B(n3252), .OUT(n3250) );
  NAND2 U1700 ( .A(n3254), .B(n3255), .OUT(n3253) );
  NOR2 U1701 ( .A(n3257), .B(n3258), .OUT(n3256) );
  NAND2 U1702 ( .A(n3260), .B(n3261), .OUT(n3259) );
  NOR2 U1703 ( .A(n3263), .B(n3264), .OUT(n3262) );
  NAND2 U1704 ( .A(n3266), .B(n3267), .OUT(n3265) );
  NOR2 U1705 ( .A(n3269), .B(n3270), .OUT(n3268) );
  NAND2 U1706 ( .A(n3272), .B(n3273), .OUT(n3271) );
  NOR2 U1707 ( .A(n3275), .B(n3276), .OUT(n3274) );
  NAND2 U1708 ( .A(n3278), .B(n3279), .OUT(n3277) );
  NOR2 U1709 ( .A(n3281), .B(n3282), .OUT(n3280) );
  NAND2 U1710 ( .A(n3284), .B(n3285), .OUT(n3283) );
  NOR2 U1711 ( .A(n3287), .B(n3288), .OUT(n3286) );
  NAND2 U1712 ( .A(n3290), .B(n3291), .OUT(n3289) );
  NOR2 U1713 ( .A(n3293), .B(n3294), .OUT(n3292) );
  NAND2 U1714 ( .A(n3296), .B(n3297), .OUT(n3295) );
  NOR2 U1715 ( .A(n3299), .B(n3300), .OUT(n3298) );
  NAND2 U1716 ( .A(n3302), .B(n3303), .OUT(n3301) );
  NOR2 U1717 ( .A(n3305), .B(n3306), .OUT(n3304) );
  NAND2 U1718 ( .A(n3308), .B(n3309), .OUT(n3307) );
  NOR2 U1719 ( .A(n3311), .B(n3312), .OUT(n3310) );
  NAND2 U1720 ( .A(n3314), .B(n3315), .OUT(n3313) );
  NOR2 U1721 ( .A(n3317), .B(n3318), .OUT(n3316) );
  NAND2 U1722 ( .A(n3320), .B(n3321), .OUT(n3319) );
  NOR2 U1723 ( .A(n3323), .B(n3324), .OUT(n3322) );
  NAND2 U1724 ( .A(n3326), .B(n3327), .OUT(n3325) );
  NOR2 U1725 ( .A(n3329), .B(n3330), .OUT(n3328) );
  NAND2 U1726 ( .A(n3332), .B(n3333), .OUT(n3331) );
  NOR2 U1727 ( .A(n3335), .B(n3336), .OUT(n3334) );
  NAND2 U1728 ( .A(n3338), .B(n3339), .OUT(n3337) );
  NOR2 U1729 ( .A(n3341), .B(n3342), .OUT(n3340) );
  NAND2 U1730 ( .A(n3344), .B(n3345), .OUT(n3343) );
  NOR2 U1731 ( .A(n3347), .B(n3348), .OUT(n3346) );
  NAND2 U1732 ( .A(n3350), .B(n3351), .OUT(n3349) );
  NOR2 U1733 ( .A(n3353), .B(n3354), .OUT(n3352) );
  NAND2 U1734 ( .A(n3356), .B(n3357), .OUT(n3355) );
  NOR2 U1735 ( .A(n3359), .B(n3360), .OUT(n3358) );
  NAND2 U1736 ( .A(n3362), .B(n3363), .OUT(n3361) );
  NOR2 U1737 ( .A(n3365), .B(n3366), .OUT(n3364) );
  NAND2 U1738 ( .A(n3368), .B(n3369), .OUT(n3367) );
  NOR2 U1739 ( .A(n3371), .B(n3372), .OUT(n3370) );
  NAND2 U1740 ( .A(n3374), .B(n3375), .OUT(n3373) );
  NOR2 U1741 ( .A(n3377), .B(n3378), .OUT(n3376) );
  NOR2 U1742 ( .A(n3380), .B(n3381), .OUT(n3379) );
  NOR2 U1743 ( .A(n3383), .B(n3384), .OUT(n3382) );
  NOR2 U1744 ( .A(n3386), .B(n3387), .OUT(n3385) );
  NOR2 U1745 ( .A(n3389), .B(n3390), .OUT(n3388) );
  NOR2 U1746 ( .A(n3392), .B(n3393), .OUT(n3391) );
  NOR2 U1747 ( .A(n3395), .B(n3396), .OUT(n3394) );
  NOR2 U1748 ( .A(n3398), .B(n3399), .OUT(n3397) );
  NOR2 U1749 ( .A(n3401), .B(n3402), .OUT(n3400) );
  NOR2 U1750 ( .A(n3404), .B(n3405), .OUT(n3403) );
  NAND2 U1751 ( .A(n3407), .B(n3408), .OUT(n3406) );
  NOR2 U1752 ( .A(n3410), .B(n3411), .OUT(n3409) );
  NOR2 U1753 ( .A(n3413), .B(n3414), .OUT(n3412) );
  NOR2 U1754 ( .A(n3416), .B(n3417), .OUT(n3415) );
  NAND2 U1755 ( .A(n3419), .B(n3420), .OUT(n3418) );
  NOR2 U1756 ( .A(n3422), .B(n3423), .OUT(n3421) );
  NOR2 U1757 ( .A(n3425), .B(n3426), .OUT(n3424) );
  NOR2 U1758 ( .A(n3428), .B(n3429), .OUT(n3427) );
  NAND2 U1759 ( .A(n3431), .B(n3432), .OUT(n3430) );
  NOR2 U1760 ( .A(n3434), .B(n3435), .OUT(n3433) );
  NOR2 U1761 ( .A(n3437), .B(n3438), .OUT(n3436) );
  NOR2 U1762 ( .A(n3440), .B(n3441), .OUT(n3439) );
  NAND2 U1763 ( .A(n3443), .B(n3444), .OUT(n3442) );
  NOR2 U1764 ( .A(n3446), .B(n3447), .OUT(n3445) );
  NOR2 U1765 ( .A(n3449), .B(n3450), .OUT(n3448) );
  NOR2 U1766 ( .A(n3452), .B(n3453), .OUT(n3451) );
  NAND2 U1767 ( .A(n3455), .B(n3456), .OUT(n3454) );
  NOR2 U1768 ( .A(n3458), .B(n3459), .OUT(n3457) );
  NOR2 U1769 ( .A(n3461), .B(n3462), .OUT(n3460) );
  NOR2 U1770 ( .A(n3464), .B(n3465), .OUT(n3463) );
  NAND2 U1771 ( .A(n3467), .B(n3468), .OUT(n3466) );
  NOR2 U1772 ( .A(n3470), .B(n3471), .OUT(n3469) );
  NOR2 U1773 ( .A(n3473), .B(n3474), .OUT(n3472) );
  NOR2 U1774 ( .A(n3476), .B(n3477), .OUT(n3475) );
  NAND2 U1775 ( .A(n3479), .B(n3480), .OUT(n3478) );
  NOR2 U1776 ( .A(n3482), .B(n3483), .OUT(n3481) );
  NOR2 U1777 ( .A(n3485), .B(n3486), .OUT(n3484) );
  NOR2 U1778 ( .A(n3488), .B(n3489), .OUT(n3487) );
  NAND2 U1779 ( .A(n3491), .B(n3492), .OUT(n3490) );
  NOR2 U1780 ( .A(n3494), .B(n3495), .OUT(n3493) );
  NOR2 U1781 ( .A(n3497), .B(n3498), .OUT(n3496) );
  NOR2 U1782 ( .A(n3500), .B(n3501), .OUT(n3499) );
  NAND2 U1783 ( .A(n3503), .B(n3504), .OUT(n3502) );
  NOR2 U1784 ( .A(n3506), .B(n3507), .OUT(n3505) );
  NOR2 U1785 ( .A(n3509), .B(n3510), .OUT(n3508) );
  NOR2 U1786 ( .A(n3512), .B(n3513), .OUT(n3511) );
  NAND2 U1787 ( .A(n3515), .B(n3516), .OUT(n3514) );
  NOR2 U1788 ( .A(n3518), .B(n3519), .OUT(n3517) );
  NAND2 U1789 ( .A(n3521), .B(n3522), .OUT(n3520) );
  NAND2 U1790 ( .A(n3523), .B(n3524), .OUT(\mult_49/A1[28] ) );
  NAND2 U1791 ( .A(n3525), .B(n3526), .OUT(\mult_49/A1[26] ) );
  NAND2 U1792 ( .A(n3527), .B(n3528), .OUT(\mult_49/A1[24] ) );
  NAND2 U1793 ( .A(n3529), .B(n3530), .OUT(\mult_49/A1[22] ) );
  NAND2 U1794 ( .A(n3531), .B(n3532), .OUT(\mult_49/A1[20] ) );
  NAND2 U1795 ( .A(n3533), .B(n3534), .OUT(\mult_49/A1[18] ) );
  NAND2 U1796 ( .A(n3535), .B(n3536), .OUT(\mult_49/A1[16] ) );
  NAND2 U1797 ( .A(n3537), .B(n3538), .OUT(\mult_49/A1[14] ) );
  NAND2 U1798 ( .A(n3539), .B(n3540), .OUT(\mult_49/A1[12] ) );
  NAND2 U1799 ( .A(n3541), .B(n3542), .OUT(\mult_49/A1[10] ) );
  NAND2 U1800 ( .A(n3543), .B(n3544), .OUT(\mult_49/A1[0] ) );
  NAND2 U1801 ( .A(n3546), .B(n3547), .OUT(n3545) );
  NAND2 U1802 ( .A(n3549), .B(n3550), .OUT(n3548) );
  NAND2 U1803 ( .A(n3552), .B(n3553), .OUT(n3551) );
  NAND2 U1804 ( .A(n3555), .B(n3556), .OUT(n3554) );
  NAND2 U1805 ( .A(n3558), .B(n3559), .OUT(n3557) );
  NAND2 U1806 ( .A(n3561), .B(n3562), .OUT(n3560) );
  NAND2 U1807 ( .A(n3564), .B(n3565), .OUT(n3563) );
  NOR2 U1808 ( .A(n3566), .B(n3567), .OUT(\gt_48/AEQB [31]) );
  NAND2 U1809 ( .A(n3569), .B(n3570), .OUT(n3568) );
  NAND2 U1810 ( .A(n3572), .B(n3573), .OUT(n3571) );
  NAND2 U1811 ( .A(n3575), .B(n3576), .OUT(n3574) );
  NAND2 U1812 ( .A(n3578), .B(n3579), .OUT(n3577) );
  NAND2 U1813 ( .A(n3581), .B(n3582), .OUT(n3580) );
  NAND2 U1814 ( .A(n3584), .B(n3585), .OUT(n3583) );
  NAND2 U1815 ( .A(n3587), .B(n3588), .OUT(n3586) );
  NAND2 U1816 ( .A(n3590), .B(n3591), .OUT(n3589) );
  NAND2 U1817 ( .A(n3593), .B(n3594), .OUT(n3592) );
  NAND2 U1818 ( .A(n3596), .B(n3597), .OUT(n3595) );
  NAND2 U1819 ( .A(n3599), .B(n3600), .OUT(n3598) );
  NAND2 U1820 ( .A(n3602), .B(n3603), .OUT(n3601) );
  NAND2 U1821 ( .A(n3605), .B(n3606), .OUT(n3604) );
  NAND2 U1822 ( .A(n3608), .B(n3609), .OUT(n3607) );
  NAND2 U1823 ( .A(n3611), .B(n3612), .OUT(n3610) );
  NAND2 U1824 ( .A(n3614), .B(n3615), .OUT(n3613) );
  NAND2 U1825 ( .A(n3617), .B(n3618), .OUT(n3616) );
  NAND2 U1826 ( .A(n3620), .B(n3621), .OUT(n3619) );
  NAND2 U1827 ( .A(n3623), .B(n3624), .OUT(n3622) );
  NAND2 U1828 ( .A(n3626), .B(n3627), .OUT(n3625) );
  NAND2 U1829 ( .A(n3629), .B(n3630), .OUT(n3628) );
  NAND2 U1830 ( .A(n3632), .B(n3633), .OUT(n3631) );
  NAND2 U1831 ( .A(n3635), .B(n3636), .OUT(n3634) );
  NAND2 U1832 ( .A(n3637), .B(n3638), .OUT(N94) );
  NAND2 U1833 ( .A(n3639), .B(n3640), .OUT(N223) );
  NAND2 U1834 ( .A(n3641), .B(n3642), .OUT(N188) );
  NAND2 U1835 ( .A(n3643), .B(n3644), .OUT(N187) );
  NAND2 U1836 ( .A(n3645), .B(n3646), .OUT(N186) );
  NAND2 U1837 ( .A(n3647), .B(n3648), .OUT(N185) );
  NAND2 U1838 ( .A(n3649), .B(n3650), .OUT(N184) );
  NAND2 U1839 ( .A(n3651), .B(n3652), .OUT(N183) );
  NAND2 U1840 ( .A(n3653), .B(n3654), .OUT(N182) );
  NAND2 U1841 ( .A(n3655), .B(n3656), .OUT(N181) );
  NAND2 U1842 ( .A(n3657), .B(n3658), .OUT(N180) );
  NAND2 U1843 ( .A(n3659), .B(n3660), .OUT(N179) );
  NAND2 U1844 ( .A(n3661), .B(n3662), .OUT(N178) );
  NAND2 U1845 ( .A(n3663), .B(n3664), .OUT(N177) );
  NAND2 U1846 ( .A(n3665), .B(n3666), .OUT(N176) );
  NAND2 U1847 ( .A(n3667), .B(n3668), .OUT(N175) );
  NAND2 U1848 ( .A(n3669), .B(n3670), .OUT(N174) );
  NAND2 U1849 ( .A(n3671), .B(n3672), .OUT(N173) );
  NAND2 U1850 ( .A(n3673), .B(n3674), .OUT(N172) );
  NAND2 U1851 ( .A(n3675), .B(n3676), .OUT(N171) );
  NAND2 U1852 ( .A(n3677), .B(n3678), .OUT(N170) );
  NAND2 U1853 ( .A(n3679), .B(n3680), .OUT(N169) );
  NAND2 U1854 ( .A(n3681), .B(n3682), .OUT(N168) );
  NAND2 U1855 ( .A(n3683), .B(n3684), .OUT(N167) );
  NAND2 U1856 ( .A(n3685), .B(n3686), .OUT(N166) );
  NAND2 U1857 ( .A(n3687), .B(n3688), .OUT(N165) );
  NAND2 U1858 ( .A(n3689), .B(n3690), .OUT(N164) );
  NAND2 U1859 ( .A(n3691), .B(n3692), .OUT(N163) );
  NAND2 U1860 ( .A(n3693), .B(n3694), .OUT(N162) );
  NAND2 U1861 ( .A(n3695), .B(n3696), .OUT(N161) );
  NAND2 U1862 ( .A(n3697), .B(n3698), .OUT(N160) );
  NAND2 U1863 ( .A(n3699), .B(n3700), .OUT(N159) );
  NAND2 U1864 ( .A(n3701), .B(n3702), .OUT(N158) );
  NAND2 U1865 ( .A(n3704), .B(n3705), .OUT(n3703) );
  NAND2 U1866 ( .A(n3707), .B(n3708), .OUT(n3706) );
  NAND2 U1867 ( .A(n3710), .B(n444), .OUT(n3709) );
  NAND2 U1868 ( .A(n3712), .B(n3713), .OUT(n3711) );
  NAND2 U1869 ( .A(n3715), .B(n412), .OUT(n3714) );
  NAND2 U1870 ( .A(n3717), .B(n448), .OUT(n3716) );
  NAND2 U1871 ( .A(n3719), .B(n3720), .OUT(n3718) );
  NAND2 U1872 ( .A(n3722), .B(n384), .OUT(n3721) );
  NAND2 U1873 ( .A(n3724), .B(n416), .OUT(n3723) );
  NAND2 U1874 ( .A(n3726), .B(n452), .OUT(n3725) );
  NAND2 U1875 ( .A(n3728), .B(n3729), .OUT(n3727) );
  NAND2 U1876 ( .A(n3731), .B(n360), .OUT(n3730) );
  NAND2 U1877 ( .A(n3733), .B(n388), .OUT(n3732) );
  NAND2 U1878 ( .A(n3735), .B(n420), .OUT(n3734) );
  NAND2 U1879 ( .A(n3737), .B(n456), .OUT(n3736) );
  NAND2 U1880 ( .A(n3739), .B(n3740), .OUT(n3738) );
  NAND2 U1881 ( .A(n3742), .B(n340), .OUT(n3741) );
  NAND2 U1882 ( .A(n3744), .B(n364), .OUT(n3743) );
  NAND2 U1883 ( .A(n3746), .B(n392), .OUT(n3745) );
  NAND2 U1884 ( .A(n3748), .B(n424), .OUT(n3747) );
  NAND2 U1885 ( .A(n3750), .B(n460), .OUT(n3749) );
  NAND2 U1886 ( .A(n3752), .B(n3753), .OUT(n3751) );
  NAND2 U1887 ( .A(n3755), .B(n324), .OUT(n3754) );
  NAND2 U1888 ( .A(n3757), .B(n344), .OUT(n3756) );
  NAND2 U1889 ( .A(n3759), .B(n368), .OUT(n3758) );
  NAND2 U1890 ( .A(n3761), .B(n396), .OUT(n3760) );
  NAND2 U1891 ( .A(n3763), .B(n428), .OUT(n3762) );
  NAND2 U1892 ( .A(n3765), .B(n464), .OUT(n3764) );
  NAND2 U1893 ( .A(n3767), .B(n3768), .OUT(n3766) );
  NAND2 U1894 ( .A(n3770), .B(n313), .OUT(n3769) );
  NAND2 U1895 ( .A(n3772), .B(n329), .OUT(n3771) );
  NAND2 U1896 ( .A(n3774), .B(n349), .OUT(n3773) );
  NAND2 U1897 ( .A(n3776), .B(n373), .OUT(n3775) );
  NAND2 U1898 ( .A(n3778), .B(n401), .OUT(n3777) );
  NAND2 U1899 ( .A(n3780), .B(n433), .OUT(n3779) );
  NAND2 U1900 ( .A(n3782), .B(n469), .OUT(n3781) );
  NAND2 U1901 ( .A(n3784), .B(n3785), .OUT(n3783) );
  NAND2 U1902 ( .A(n3787), .B(n524), .OUT(n3786) );
  NAND2 U1903 ( .A(n3789), .B(n528), .OUT(n3788) );
  NAND2 U1904 ( .A(n3791), .B(n532), .OUT(n3790) );
  NAND2 U1905 ( .A(n3793), .B(n536), .OUT(n3792) );
  NAND2 U1906 ( .A(n3795), .B(n540), .OUT(n3794) );
  NAND2 U1907 ( .A(n3797), .B(n544), .OUT(n3796) );
  NAND2 U1908 ( .A(n3799), .B(n512), .OUT(n3798) );
  NAND2 U1909 ( .A(n3801), .B(n1880), .OUT(n3800) );
  NAND2 U1910 ( .A(n3803), .B(n1956), .OUT(n3802) );
  NAND2 U1911 ( .A(n3805), .B(n509), .OUT(n3804) );
  NAND2 U1912 ( .A(n3807), .B(n504), .OUT(n3806) );
  NAND2 U1913 ( .A(n3809), .B(n500), .OUT(n3808) );
  NAND2 U1914 ( .A(n3811), .B(n496), .OUT(n3810) );
  NAND2 U1915 ( .A(n3813), .B(n492), .OUT(n3812) );
  NAND2 U1916 ( .A(n3815), .B(n488), .OUT(n3814) );
  NAND2 U1917 ( .A(n3817), .B(n484), .OUT(n3816) );
  NAND2 U1918 ( .A(n3819), .B(n3820), .OUT(n3818) );
  NAND2 U1919 ( .A(n3822), .B(n560), .OUT(n3821) );
  NAND2 U1920 ( .A(n3824), .B(n564), .OUT(n3823) );
  NAND2 U1921 ( .A(n3826), .B(n568), .OUT(n3825) );
  NAND2 U1922 ( .A(n3828), .B(n572), .OUT(n3827) );
  NAND2 U1923 ( .A(n3830), .B(n576), .OUT(n3829) );
  NAND2 U1924 ( .A(n3832), .B(n580), .OUT(n3831) );
  NAND2 U1925 ( .A(n3834), .B(n584), .OUT(n3833) );
  NAND2 U1926 ( .A(n3836), .B(n3837), .OUT(n3835) );
  NAND2 U1927 ( .A(n3839), .B(n600), .OUT(n3838) );
  NAND2 U1928 ( .A(n3841), .B(n604), .OUT(n3840) );
  NAND2 U1929 ( .A(n3843), .B(n608), .OUT(n3842) );
  NAND2 U1930 ( .A(n3845), .B(n612), .OUT(n3844) );
  NAND2 U1931 ( .A(n3847), .B(n616), .OUT(n3846) );
  NAND2 U1932 ( .A(n3849), .B(n620), .OUT(n3848) );
  NAND2 U1933 ( .A(n3851), .B(n624), .OUT(n3850) );
  NAND2 U1934 ( .A(n3853), .B(n628), .OUT(n3852) );
  NAND2 U1935 ( .A(n3855), .B(n3856), .OUT(n3854) );
  NAND2 U1936 ( .A(n3858), .B(n644), .OUT(n3857) );
  NAND2 U1937 ( .A(n3860), .B(n648), .OUT(n3859) );
  NAND2 U1938 ( .A(n3862), .B(n652), .OUT(n3861) );
  NAND2 U1939 ( .A(n3864), .B(n656), .OUT(n3863) );
  NAND2 U1940 ( .A(n3866), .B(n660), .OUT(n3865) );
  NAND2 U1941 ( .A(n3868), .B(n664), .OUT(n3867) );
  NAND2 U1942 ( .A(n3870), .B(n668), .OUT(n3869) );
  NAND2 U1943 ( .A(n3872), .B(n672), .OUT(n3871) );
  NAND2 U1944 ( .A(n3874), .B(n676), .OUT(n3873) );
  NAND2 U1945 ( .A(n3876), .B(n3877), .OUT(n3875) );
  NAND2 U1946 ( .A(n3879), .B(n692), .OUT(n3878) );
  NAND2 U1947 ( .A(n3881), .B(n696), .OUT(n3880) );
  NAND2 U1948 ( .A(n3883), .B(n700), .OUT(n3882) );
  NAND2 U1949 ( .A(n3885), .B(n704), .OUT(n3884) );
  NAND2 U1950 ( .A(n3887), .B(n708), .OUT(n3886) );
  NAND2 U1951 ( .A(n3889), .B(n712), .OUT(n3888) );
  NAND2 U1952 ( .A(n3891), .B(n716), .OUT(n3890) );
  NAND2 U1953 ( .A(n3893), .B(n720), .OUT(n3892) );
  NAND2 U1954 ( .A(n3895), .B(n724), .OUT(n3894) );
  NAND2 U1955 ( .A(n3897), .B(n728), .OUT(n3896) );
  NAND2 U1956 ( .A(n3899), .B(n3900), .OUT(n3898) );
  NAND2 U1957 ( .A(n3902), .B(n744), .OUT(n3901) );
  NAND2 U1958 ( .A(n3904), .B(n748), .OUT(n3903) );
  NAND2 U1959 ( .A(n3906), .B(n752), .OUT(n3905) );
  NAND2 U1960 ( .A(n3908), .B(n756), .OUT(n3907) );
  NAND2 U1961 ( .A(n3910), .B(n760), .OUT(n3909) );
  NAND2 U1962 ( .A(n3912), .B(n764), .OUT(n3911) );
  NAND2 U1963 ( .A(n3914), .B(n768), .OUT(n3913) );
  NAND2 U1964 ( .A(n3916), .B(n772), .OUT(n3915) );
  NAND2 U1965 ( .A(n3918), .B(n776), .OUT(n3917) );
  NAND2 U1966 ( .A(n3920), .B(n780), .OUT(n3919) );
  NAND2 U1967 ( .A(n3922), .B(n784), .OUT(n3921) );
  NAND2 U1968 ( .A(n3924), .B(n3925), .OUT(n3923) );
  NAND2 U1969 ( .A(n3927), .B(n800), .OUT(n3926) );
  NAND2 U1970 ( .A(n3929), .B(n804), .OUT(n3928) );
  NAND2 U1971 ( .A(n3931), .B(n808), .OUT(n3930) );
  NAND2 U1972 ( .A(n3933), .B(n812), .OUT(n3932) );
  NAND2 U1973 ( .A(n3935), .B(n816), .OUT(n3934) );
  NAND2 U1974 ( .A(n3937), .B(n820), .OUT(n3936) );
  NAND2 U1975 ( .A(n3939), .B(n824), .OUT(n3938) );
  NAND2 U1976 ( .A(n3941), .B(n828), .OUT(n3940) );
  NAND2 U1977 ( .A(n3943), .B(n832), .OUT(n3942) );
  NAND2 U1978 ( .A(n3945), .B(n836), .OUT(n3944) );
  NAND2 U1979 ( .A(n3947), .B(n840), .OUT(n3946) );
  NAND2 U1980 ( .A(n3949), .B(n844), .OUT(n3948) );
  NAND2 U1981 ( .A(n3951), .B(n3952), .OUT(n3950) );
  NAND2 U1982 ( .A(n3954), .B(n860), .OUT(n3953) );
  NAND2 U1983 ( .A(n3956), .B(n864), .OUT(n3955) );
  NAND2 U1984 ( .A(n3958), .B(n868), .OUT(n3957) );
  NAND2 U1985 ( .A(n3960), .B(n872), .OUT(n3959) );
  NAND2 U1986 ( .A(n3962), .B(n876), .OUT(n3961) );
  NAND2 U1987 ( .A(n3964), .B(n880), .OUT(n3963) );
  NAND2 U1988 ( .A(n3966), .B(n884), .OUT(n3965) );
  NAND2 U1989 ( .A(n3968), .B(n888), .OUT(n3967) );
  NAND2 U1990 ( .A(n3970), .B(n892), .OUT(n3969) );
  NAND2 U1991 ( .A(n3972), .B(n896), .OUT(n3971) );
  NAND2 U1992 ( .A(n3974), .B(n900), .OUT(n3973) );
  NAND2 U1993 ( .A(n3976), .B(n904), .OUT(n3975) );
  NAND2 U1994 ( .A(n3978), .B(n908), .OUT(n3977) );
  NAND2 U1995 ( .A(n3980), .B(n3981), .OUT(n3979) );
  NAND2 U1996 ( .A(n3983), .B(n924), .OUT(n3982) );
  NAND2 U1997 ( .A(n3985), .B(n928), .OUT(n3984) );
  NAND2 U1998 ( .A(n3987), .B(n932), .OUT(n3986) );
  NAND2 U1999 ( .A(n3989), .B(n936), .OUT(n3988) );
  NAND2 U2000 ( .A(n3991), .B(n940), .OUT(n3990) );
  NAND2 U2001 ( .A(n3993), .B(n944), .OUT(n3992) );
  NAND2 U2002 ( .A(n3995), .B(n948), .OUT(n3994) );
  NAND2 U2003 ( .A(n3997), .B(n952), .OUT(n3996) );
  NAND2 U2004 ( .A(n3999), .B(n956), .OUT(n3998) );
  NAND2 U2005 ( .A(n4001), .B(n960), .OUT(n4000) );
  NAND2 U2006 ( .A(n4003), .B(n964), .OUT(n4002) );
  NAND2 U2007 ( .A(n4005), .B(n968), .OUT(n4004) );
  NAND2 U2008 ( .A(n4007), .B(n972), .OUT(n4006) );
  NAND2 U2009 ( .A(n4009), .B(n976), .OUT(n4008) );
  NAND2 U2010 ( .A(n4011), .B(n4012), .OUT(n4010) );
  NAND2 U2011 ( .A(n4014), .B(n992), .OUT(n4013) );
  NAND2 U2012 ( .A(n4016), .B(n996), .OUT(n4015) );
  NAND2 U2013 ( .A(n4018), .B(n1000), .OUT(n4017) );
  NAND2 U2014 ( .A(n4020), .B(n1004), .OUT(n4019) );
  NAND2 U2015 ( .A(n4022), .B(n1008), .OUT(n4021) );
  NAND2 U2016 ( .A(n4024), .B(n1012), .OUT(n4023) );
  NAND2 U2017 ( .A(n4026), .B(n1016), .OUT(n4025) );
  NAND2 U2018 ( .A(n4028), .B(n1020), .OUT(n4027) );
  NAND2 U2019 ( .A(n4030), .B(n1024), .OUT(n4029) );
  NAND2 U2020 ( .A(n4032), .B(n1028), .OUT(n4031) );
  NAND2 U2021 ( .A(n4034), .B(n1032), .OUT(n4033) );
  NAND2 U2022 ( .A(n4036), .B(n1036), .OUT(n4035) );
  NAND2 U2023 ( .A(n4038), .B(n1040), .OUT(n4037) );
  NAND2 U2024 ( .A(n4040), .B(n1044), .OUT(n4039) );
  NAND2 U2025 ( .A(n4042), .B(n1048), .OUT(n4041) );
  NAND2 U2026 ( .A(n4044), .B(n4045), .OUT(n4043) );
  NAND2 U2027 ( .A(n4047), .B(n1064), .OUT(n4046) );
  NAND2 U2028 ( .A(n4049), .B(n1068), .OUT(n4048) );
  NAND2 U2029 ( .A(n4051), .B(n1072), .OUT(n4050) );
  NAND2 U2030 ( .A(n4053), .B(n1076), .OUT(n4052) );
  NAND2 U2031 ( .A(n4055), .B(n1080), .OUT(n4054) );
  NAND2 U2032 ( .A(n4057), .B(n1084), .OUT(n4056) );
  NAND2 U2033 ( .A(n4059), .B(n1088), .OUT(n4058) );
  NAND2 U2034 ( .A(n4061), .B(n1092), .OUT(n4060) );
  NAND2 U2035 ( .A(n4063), .B(n1096), .OUT(n4062) );
  NAND2 U2036 ( .A(n4065), .B(n1100), .OUT(n4064) );
  NAND2 U2037 ( .A(n4067), .B(n1104), .OUT(n4066) );
  NAND2 U2038 ( .A(n4069), .B(n1108), .OUT(n4068) );
  NAND2 U2039 ( .A(n4071), .B(n1112), .OUT(n4070) );
  NAND2 U2040 ( .A(n4073), .B(n1116), .OUT(n4072) );
  NAND2 U2041 ( .A(n4075), .B(n1120), .OUT(n4074) );
  NAND2 U2042 ( .A(n4077), .B(n1124), .OUT(n4076) );
  NAND2 U2043 ( .A(n4079), .B(n4080), .OUT(n4078) );
  NAND2 U2044 ( .A(n4082), .B(n1140), .OUT(n4081) );
  NAND2 U2045 ( .A(n4084), .B(n1144), .OUT(n4083) );
  NAND2 U2046 ( .A(n4086), .B(n1148), .OUT(n4085) );
  NAND2 U2047 ( .A(n4088), .B(n1152), .OUT(n4087) );
  NAND2 U2048 ( .A(n4090), .B(n1156), .OUT(n4089) );
  NAND2 U2049 ( .A(n4092), .B(n1160), .OUT(n4091) );
  NAND2 U2050 ( .A(n4094), .B(n1164), .OUT(n4093) );
  NAND2 U2051 ( .A(n4096), .B(n1168), .OUT(n4095) );
  NAND2 U2052 ( .A(n4098), .B(n1172), .OUT(n4097) );
  NAND2 U2053 ( .A(n4100), .B(n1176), .OUT(n4099) );
  NAND2 U2054 ( .A(n4102), .B(n1180), .OUT(n4101) );
  NAND2 U2055 ( .A(n4104), .B(n1184), .OUT(n4103) );
  NAND2 U2056 ( .A(n4106), .B(n1188), .OUT(n4105) );
  NAND2 U2057 ( .A(n4108), .B(n1192), .OUT(n4107) );
  NAND2 U2058 ( .A(n4110), .B(n1196), .OUT(n4109) );
  NAND2 U2059 ( .A(n4112), .B(n1200), .OUT(n4111) );
  NAND2 U2060 ( .A(n4114), .B(n1204), .OUT(n4113) );
  NAND2 U2061 ( .A(n4116), .B(n4117), .OUT(n4115) );
  NAND2 U2062 ( .A(n4119), .B(n1220), .OUT(n4118) );
  NAND2 U2063 ( .A(n4121), .B(n1224), .OUT(n4120) );
  NAND2 U2064 ( .A(n4123), .B(n1228), .OUT(n4122) );
  NAND2 U2065 ( .A(n4125), .B(n1232), .OUT(n4124) );
  NAND2 U2066 ( .A(n4127), .B(n1236), .OUT(n4126) );
  NAND2 U2067 ( .A(n4129), .B(n1240), .OUT(n4128) );
  NAND2 U2068 ( .A(n4131), .B(n1244), .OUT(n4130) );
  NAND2 U2069 ( .A(n4133), .B(n1248), .OUT(n4132) );
  NAND2 U2070 ( .A(n4135), .B(n1252), .OUT(n4134) );
  NAND2 U2071 ( .A(n4137), .B(n1256), .OUT(n4136) );
  NAND2 U2072 ( .A(n4139), .B(n1260), .OUT(n4138) );
  NAND2 U2073 ( .A(n4141), .B(n1264), .OUT(n4140) );
  NAND2 U2074 ( .A(n4143), .B(n1268), .OUT(n4142) );
  NAND2 U2075 ( .A(n4145), .B(n1272), .OUT(n4144) );
  NAND2 U2076 ( .A(n4147), .B(n1276), .OUT(n4146) );
  NAND2 U2077 ( .A(n4149), .B(n1280), .OUT(n4148) );
  NAND2 U2078 ( .A(n4151), .B(n1284), .OUT(n4150) );
  NAND2 U2079 ( .A(n4153), .B(n1288), .OUT(n4152) );
  NAND2 U2080 ( .A(n4155), .B(n4156), .OUT(n4154) );
  NAND2 U2081 ( .A(n4158), .B(n1304), .OUT(n4157) );
  NAND2 U2082 ( .A(n4160), .B(n1308), .OUT(n4159) );
  NAND2 U2083 ( .A(n4162), .B(n1312), .OUT(n4161) );
  NAND2 U2084 ( .A(n4164), .B(n1316), .OUT(n4163) );
  NAND2 U2085 ( .A(n4166), .B(n1320), .OUT(n4165) );
  NAND2 U2086 ( .A(n4168), .B(n1324), .OUT(n4167) );
  NAND2 U2087 ( .A(n4170), .B(n1328), .OUT(n4169) );
  NAND2 U2088 ( .A(n4172), .B(n1332), .OUT(n4171) );
  NAND2 U2089 ( .A(n4174), .B(n1336), .OUT(n4173) );
  NAND2 U2090 ( .A(n4176), .B(n1340), .OUT(n4175) );
  NAND2 U2091 ( .A(n4178), .B(n1344), .OUT(n4177) );
  NAND2 U2092 ( .A(n4180), .B(n1348), .OUT(n4179) );
  NAND2 U2093 ( .A(n4182), .B(n1352), .OUT(n4181) );
  NAND2 U2094 ( .A(n4184), .B(n1356), .OUT(n4183) );
  NAND2 U2095 ( .A(n4186), .B(n1360), .OUT(n4185) );
  NAND2 U2096 ( .A(n4188), .B(n1364), .OUT(n4187) );
  NAND2 U2097 ( .A(n4190), .B(n1368), .OUT(n4189) );
  NAND2 U2098 ( .A(n4192), .B(n1372), .OUT(n4191) );
  NAND2 U2099 ( .A(n4194), .B(n1376), .OUT(n4193) );
  NAND2 U2100 ( .A(n4196), .B(n4197), .OUT(n4195) );
  NAND2 U2101 ( .A(n4199), .B(n1392), .OUT(n4198) );
  NAND2 U2102 ( .A(n4201), .B(n1396), .OUT(n4200) );
  NAND2 U2103 ( .A(n4203), .B(n1400), .OUT(n4202) );
  NAND2 U2104 ( .A(n4205), .B(n1404), .OUT(n4204) );
  NAND2 U2105 ( .A(n4207), .B(n1408), .OUT(n4206) );
  NAND2 U2106 ( .A(n4209), .B(n1412), .OUT(n4208) );
  NAND2 U2107 ( .A(n4211), .B(n1416), .OUT(n4210) );
  NAND2 U2108 ( .A(n4213), .B(n1420), .OUT(n4212) );
  NAND2 U2109 ( .A(n4215), .B(n1424), .OUT(n4214) );
  NAND2 U2110 ( .A(n4217), .B(n1428), .OUT(n4216) );
  NAND2 U2111 ( .A(n4219), .B(n1432), .OUT(n4218) );
  NAND2 U2112 ( .A(n4221), .B(n1436), .OUT(n4220) );
  NAND2 U2113 ( .A(n4223), .B(n1440), .OUT(n4222) );
  NAND2 U2114 ( .A(n4225), .B(n1444), .OUT(n4224) );
  NAND2 U2115 ( .A(n4227), .B(n1448), .OUT(n4226) );
  NAND2 U2116 ( .A(n4229), .B(n1452), .OUT(n4228) );
  NAND2 U2117 ( .A(n4231), .B(n1456), .OUT(n4230) );
  NAND2 U2118 ( .A(n4233), .B(n1460), .OUT(n4232) );
  NAND2 U2119 ( .A(n4235), .B(n1464), .OUT(n4234) );
  NAND2 U2120 ( .A(n4237), .B(n1468), .OUT(n4236) );
  NAND2 U2121 ( .A(n4239), .B(n4240), .OUT(n4238) );
  NAND2 U2122 ( .A(n4242), .B(n1484), .OUT(n4241) );
  NAND2 U2123 ( .A(n4244), .B(n1488), .OUT(n4243) );
  NAND2 U2124 ( .A(n4246), .B(n1492), .OUT(n4245) );
  NAND2 U2125 ( .A(n4248), .B(n1496), .OUT(n4247) );
  NAND2 U2126 ( .A(n4250), .B(n1500), .OUT(n4249) );
  NAND2 U2127 ( .A(n4252), .B(n1504), .OUT(n4251) );
  NAND2 U2128 ( .A(n4254), .B(n1508), .OUT(n4253) );
  NAND2 U2129 ( .A(n4256), .B(n1512), .OUT(n4255) );
  NAND2 U2130 ( .A(n4258), .B(n1516), .OUT(n4257) );
  NAND2 U2131 ( .A(n4260), .B(n1520), .OUT(n4259) );
  NAND2 U2132 ( .A(n4262), .B(n1524), .OUT(n4261) );
  NAND2 U2133 ( .A(n4264), .B(n1528), .OUT(n4263) );
  NAND2 U2134 ( .A(n4266), .B(n1532), .OUT(n4265) );
  NAND2 U2135 ( .A(n4268), .B(n1536), .OUT(n4267) );
  NAND2 U2136 ( .A(n4270), .B(n1540), .OUT(n4269) );
  NAND2 U2137 ( .A(n4272), .B(n1544), .OUT(n4271) );
  NAND2 U2138 ( .A(n4274), .B(n1548), .OUT(n4273) );
  NAND2 U2139 ( .A(n4276), .B(n1552), .OUT(n4275) );
  NAND2 U2140 ( .A(n4278), .B(n1556), .OUT(n4277) );
  NAND2 U2141 ( .A(n4280), .B(n1560), .OUT(n4279) );
  NAND2 U2142 ( .A(n4282), .B(n1564), .OUT(n4281) );
  NAND2 U2143 ( .A(n4284), .B(n4285), .OUT(n4283) );
  NAND2 U2144 ( .A(n4287), .B(n1580), .OUT(n4286) );
  NAND2 U2145 ( .A(n4289), .B(n1584), .OUT(n4288) );
  NAND2 U2146 ( .A(n4291), .B(n1588), .OUT(n4290) );
  NAND2 U2147 ( .A(n4293), .B(n1592), .OUT(n4292) );
  NAND2 U2148 ( .A(n4295), .B(n1596), .OUT(n4294) );
  NAND2 U2149 ( .A(n4297), .B(n1600), .OUT(n4296) );
  NAND2 U2150 ( .A(n4299), .B(n1604), .OUT(n4298) );
  NAND2 U2151 ( .A(n4301), .B(n1608), .OUT(n4300) );
  NAND2 U2152 ( .A(n4303), .B(n1612), .OUT(n4302) );
  NAND2 U2153 ( .A(n4305), .B(n1616), .OUT(n4304) );
  NAND2 U2154 ( .A(n4307), .B(n1620), .OUT(n4306) );
  NAND2 U2155 ( .A(n4309), .B(n1624), .OUT(n4308) );
  NAND2 U2156 ( .A(n4311), .B(n1628), .OUT(n4310) );
  NAND2 U2157 ( .A(n4313), .B(n1632), .OUT(n4312) );
  NAND2 U2158 ( .A(n4315), .B(n1636), .OUT(n4314) );
  NAND2 U2159 ( .A(n4317), .B(n1640), .OUT(n4316) );
  NAND2 U2160 ( .A(n4319), .B(n1644), .OUT(n4318) );
  NAND2 U2161 ( .A(n4321), .B(n1648), .OUT(n4320) );
  NAND2 U2162 ( .A(n4323), .B(n1652), .OUT(n4322) );
  NAND2 U2163 ( .A(n4325), .B(n1656), .OUT(n4324) );
  NAND2 U2164 ( .A(n4327), .B(n1660), .OUT(n4326) );
  NAND2 U2165 ( .A(n4329), .B(n1664), .OUT(n4328) );
  NAND2 U2166 ( .A(n4331), .B(n4332), .OUT(n4330) );
  NAND2 U2167 ( .A(n4334), .B(n1680), .OUT(n4333) );
  NAND2 U2168 ( .A(n4336), .B(n1684), .OUT(n4335) );
  NAND2 U2169 ( .A(n4338), .B(n1688), .OUT(n4337) );
  NAND2 U2170 ( .A(n4340), .B(n1692), .OUT(n4339) );
  NAND2 U2171 ( .A(n4342), .B(n1696), .OUT(n4341) );
  NAND2 U2172 ( .A(n4344), .B(n1700), .OUT(n4343) );
  NAND2 U2173 ( .A(n4346), .B(n1704), .OUT(n4345) );
  NAND2 U2174 ( .A(n4348), .B(n1708), .OUT(n4347) );
  NAND2 U2175 ( .A(n4350), .B(n1712), .OUT(n4349) );
  NAND2 U2176 ( .A(n4352), .B(n1716), .OUT(n4351) );
  NAND2 U2177 ( .A(n4354), .B(n1720), .OUT(n4353) );
  NAND2 U2178 ( .A(n4356), .B(n1724), .OUT(n4355) );
  NAND2 U2179 ( .A(n4358), .B(n1728), .OUT(n4357) );
  NAND2 U2180 ( .A(n4360), .B(n1732), .OUT(n4359) );
  NAND2 U2181 ( .A(n4362), .B(n1736), .OUT(n4361) );
  NAND2 U2182 ( .A(n4364), .B(n1740), .OUT(n4363) );
  NAND2 U2183 ( .A(n4366), .B(n1744), .OUT(n4365) );
  NAND2 U2184 ( .A(n4368), .B(n1748), .OUT(n4367) );
  NAND2 U2185 ( .A(n4370), .B(n1752), .OUT(n4369) );
  NAND2 U2186 ( .A(n4372), .B(n1756), .OUT(n4371) );
  NAND2 U2187 ( .A(n4374), .B(n1760), .OUT(n4373) );
  NAND2 U2188 ( .A(n4376), .B(n1764), .OUT(n4375) );
  NAND2 U2189 ( .A(n4378), .B(n1768), .OUT(n4377) );
  NAND2 U2190 ( .A(n4380), .B(n4381), .OUT(n4379) );
  NAND2 U2191 ( .A(n4383), .B(n1784), .OUT(n4382) );
  NAND2 U2192 ( .A(n4385), .B(n1788), .OUT(n4384) );
  NAND2 U2193 ( .A(n4387), .B(n1792), .OUT(n4386) );
  NAND2 U2194 ( .A(n4389), .B(n1796), .OUT(n4388) );
  NAND2 U2195 ( .A(n4391), .B(n1800), .OUT(n4390) );
  NAND2 U2196 ( .A(n4393), .B(n1804), .OUT(n4392) );
  NAND2 U2197 ( .A(n4395), .B(n1808), .OUT(n4394) );
  NAND2 U2198 ( .A(n4397), .B(n1812), .OUT(n4396) );
  NAND2 U2199 ( .A(n4399), .B(n1816), .OUT(n4398) );
  NAND2 U2200 ( .A(n4401), .B(n1820), .OUT(n4400) );
  NAND2 U2201 ( .A(n4403), .B(n1824), .OUT(n4402) );
  NAND2 U2202 ( .A(n4405), .B(n1828), .OUT(n4404) );
  NAND2 U2203 ( .A(n4407), .B(n1832), .OUT(n4406) );
  NAND2 U2204 ( .A(n4409), .B(n1836), .OUT(n4408) );
  NAND2 U2205 ( .A(n4411), .B(n1840), .OUT(n4410) );
  NAND2 U2206 ( .A(n4413), .B(n1844), .OUT(n4412) );
  NAND2 U2207 ( .A(n4415), .B(n1848), .OUT(n4414) );
  NAND2 U2208 ( .A(n4417), .B(n1852), .OUT(n4416) );
  NAND2 U2209 ( .A(n4419), .B(n1856), .OUT(n4418) );
  NAND2 U2210 ( .A(n4421), .B(n1860), .OUT(n4420) );
  NAND2 U2211 ( .A(n4423), .B(n1864), .OUT(n4422) );
  NAND2 U2212 ( .A(n4425), .B(n1868), .OUT(n4424) );
  NAND2 U2213 ( .A(n4427), .B(n1872), .OUT(n4426) );
  NAND2 U2214 ( .A(n4429), .B(n1876), .OUT(n4428) );
  NAND2 U2215 ( .A(n4431), .B(n4432), .OUT(n4430) );
  NAND2 U2216 ( .A(n4434), .B(n4435), .OUT(n4433) );
  NAND2 U2217 ( .A(n4437), .B(n4438), .OUT(n4436) );
  NAND2 U2218 ( .A(n4440), .B(n4441), .OUT(n4439) );
  NAND2 U2219 ( .A(n4443), .B(n4444), .OUT(n4442) );
  NAND2 U2220 ( .A(n4446), .B(n4447), .OUT(n4445) );
  NAND2 U2221 ( .A(n4449), .B(n4450), .OUT(n4448) );
  NAND2 U2222 ( .A(n4452), .B(n4453), .OUT(n4451) );
  NAND2 U2223 ( .A(n4455), .B(n4456), .OUT(n4454) );
  NAND2 U2224 ( .A(n4458), .B(n4459), .OUT(n4457) );
  NAND2 U2225 ( .A(n4461), .B(n4462), .OUT(n4460) );
  NAND2 U2226 ( .A(n4464), .B(n4465), .OUT(n4463) );
  NAND2 U2227 ( .A(n4467), .B(n4468), .OUT(n4466) );
  NAND2 U2228 ( .A(n4470), .B(n4471), .OUT(n4469) );
  NAND2 U2229 ( .A(n4473), .B(n4474), .OUT(n4472) );
  NAND2 U2230 ( .A(n4476), .B(n4477), .OUT(n4475) );
  NAND2 U2231 ( .A(n4479), .B(n4480), .OUT(n4478) );
  NAND2 U2232 ( .A(n4482), .B(n4483), .OUT(n4481) );
  NAND2 U2233 ( .A(n4485), .B(n4486), .OUT(n4484) );
  NAND2 U2234 ( .A(n4488), .B(n4489), .OUT(n4487) );
  NAND2 U2235 ( .A(n4491), .B(n4492), .OUT(n4490) );
  NAND2 U2236 ( .A(n4494), .B(n4495), .OUT(n4493) );
  NAND2 U2237 ( .A(n4497), .B(n4498), .OUT(n4496) );
  NAND2 U2238 ( .A(n4500), .B(n4501), .OUT(n4499) );
  NAND2 U2239 ( .A(n4503), .B(n4504), .OUT(n4502) );
  NAND2 U2240 ( .A(n4506), .B(n4507), .OUT(n4505) );
  NAND2 U2241 ( .A(n4509), .B(n548), .OUT(n4508) );
  NAND2 U2242 ( .A(n4511), .B(n588), .OUT(n4510) );
  NAND2 U2243 ( .A(n4513), .B(n632), .OUT(n4512) );
  NAND2 U2244 ( .A(n4515), .B(n680), .OUT(n4514) );
  NAND2 U2245 ( .A(n4517), .B(n732), .OUT(n4516) );
  NAND2 U2246 ( .A(n4519), .B(n788), .OUT(n4518) );
  NAND2 U2247 ( .A(n4521), .B(n848), .OUT(n4520) );
  NAND2 U2248 ( .A(n4523), .B(n912), .OUT(n4522) );
  NAND2 U2249 ( .A(n4525), .B(n980), .OUT(n4524) );
  NAND2 U2250 ( .A(n4527), .B(n1052), .OUT(n4526) );
  NAND2 U2251 ( .A(n4529), .B(n1128), .OUT(n4528) );
  NAND2 U2252 ( .A(n4531), .B(n1208), .OUT(n4530) );
  NAND2 U2253 ( .A(n4533), .B(n1292), .OUT(n4532) );
  NAND2 U2254 ( .A(n4535), .B(n1380), .OUT(n4534) );
  NAND2 U2255 ( .A(n4537), .B(n1472), .OUT(n4536) );
  NAND2 U2256 ( .A(n4539), .B(n1568), .OUT(n4538) );
  NAND2 U2257 ( .A(n4541), .B(n1668), .OUT(n4540) );
  NAND2 U2258 ( .A(n4543), .B(n1772), .OUT(n4542) );
  NAND2 U2259 ( .A(n4545), .B(n4546), .OUT(n4544) );
  NAND2 U2260 ( .A(n4548), .B(n1884), .OUT(n4547) );
  NAND2 U2261 ( .A(n4550), .B(n1888), .OUT(n4549) );
  NAND2 U2262 ( .A(n4552), .B(n1892), .OUT(n4551) );
  NAND2 U2263 ( .A(n4554), .B(n1896), .OUT(n4553) );
  NAND2 U2264 ( .A(n4556), .B(n1900), .OUT(n4555) );
  NAND2 U2265 ( .A(n4558), .B(n1904), .OUT(n4557) );
  NAND2 U2266 ( .A(n4560), .B(n1908), .OUT(n4559) );
  NAND2 U2267 ( .A(n4562), .B(n1912), .OUT(n4561) );
  NAND2 U2268 ( .A(n4564), .B(n1916), .OUT(n4563) );
  NAND2 U2269 ( .A(n4566), .B(n1920), .OUT(n4565) );
  NAND2 U2270 ( .A(n4568), .B(n1924), .OUT(n4567) );
  NAND2 U2271 ( .A(n4570), .B(n1928), .OUT(n4569) );
  NAND2 U2272 ( .A(n4572), .B(n1932), .OUT(n4571) );
  NAND2 U2273 ( .A(n4574), .B(n1936), .OUT(n4573) );
  NAND2 U2274 ( .A(n4576), .B(n1940), .OUT(n4575) );
  NAND2 U2275 ( .A(n4578), .B(n1944), .OUT(n4577) );
  NAND2 U2276 ( .A(n4580), .B(n1948), .OUT(n4579) );
  NAND2 U2277 ( .A(n4582), .B(n1952), .OUT(n4581) );
  NAND2 U2278 ( .A(n4584), .B(n4585), .OUT(n4583) );
  NOR2 U2279 ( .A(n4587), .B(n4588), .OUT(n4586) );
  NOR2 U2280 ( .A(n4590), .B(n4591), .OUT(n4589) );
  NOR2 U2281 ( .A(n4593), .B(n4594), .OUT(n4592) );
  NOR2 U2282 ( .A(n4596), .B(n4597), .OUT(n4595) );
  NOR2 U2283 ( .A(n4599), .B(n4600), .OUT(n4598) );
  NOR2 U2284 ( .A(n4602), .B(n4603), .OUT(n4601) );
  NOR2 U2285 ( .A(n4605), .B(n4606), .OUT(n4604) );
  NOR2 U2286 ( .A(n4608), .B(n4609), .OUT(n4607) );
  NOR2 U2287 ( .A(n4611), .B(n4612), .OUT(n4610) );
  NOR2 U2288 ( .A(n4614), .B(n4615), .OUT(n4613) );
  NOR2 U2289 ( .A(n4617), .B(n4618), .OUT(n4616) );
  NOR2 U2290 ( .A(n4620), .B(n4621), .OUT(n4619) );
  NOR2 U2291 ( .A(n4623), .B(n4624), .OUT(n4622) );
  NOR2 U2292 ( .A(n4626), .B(n4627), .OUT(n4625) );
  NOR2 U2293 ( .A(n4629), .B(n4630), .OUT(n4628) );
  NOR2 U2294 ( .A(n4632), .B(n4633), .OUT(n4631) );
  NOR2 U2295 ( .A(n4635), .B(n4636), .OUT(n4634) );
  NOR2 U2296 ( .A(n4638), .B(n4639), .OUT(n4637) );
  NOR2 U2297 ( .A(n4641), .B(n4642), .OUT(n4640) );
  NOR2 U2298 ( .A(n4644), .B(n4645), .OUT(n4643) );
  NOR2 U2299 ( .A(n4647), .B(n4648), .OUT(n4646) );
  NOR2 U2300 ( .A(n4650), .B(n4651), .OUT(n4649) );
  NOR2 U2301 ( .A(n4653), .B(n4654), .OUT(n4652) );
  NOR2 U2302 ( .A(n4656), .B(n4657), .OUT(n4655) );
  NOR2 U2303 ( .A(n4659), .B(n4660), .OUT(n4658) );
  NOR2 U2304 ( .A(n4662), .B(n4663), .OUT(n4661) );
  NOR2 U2305 ( .A(n4665), .B(n4666), .OUT(n4664) );
  NOR2 U2306 ( .A(n4668), .B(n4669), .OUT(n4667) );
  NOR2 U2307 ( .A(n4671), .B(n4672), .OUT(n4670) );
  NOR2 U2308 ( .A(n4674), .B(n4675), .OUT(n4673) );
  NOR2 U2309 ( .A(n4677), .B(n4678), .OUT(n4676) );
  NOR2 U2310 ( .A(n4680), .B(n4681), .OUT(n4679) );
  NOR2 U2311 ( .A(n4683), .B(n4684), .OUT(n4682) );
  NOR2 U2312 ( .A(n4686), .B(n4687), .OUT(n4685) );
  NOR2 U2313 ( .A(n4689), .B(n4690), .OUT(n4688) );
  NOR2 U2314 ( .A(n4692), .B(n4693), .OUT(n4691) );
  NOR2 U2315 ( .A(n4695), .B(n4696), .OUT(n4694) );
  NOR2 U2316 ( .A(n4698), .B(n4699), .OUT(n4697) );
  NOR2 U2317 ( .A(n4701), .B(n4702), .OUT(n4700) );
  NOR2 U2318 ( .A(n4704), .B(n4705), .OUT(n4703) );
  NOR2 U2319 ( .A(n4707), .B(n4708), .OUT(n4706) );
  NOR2 U2320 ( .A(n4710), .B(n4711), .OUT(n4709) );
  NOR2 U2321 ( .A(n4713), .B(n4714), .OUT(n4712) );
  NOR2 U2322 ( .A(n4716), .B(n4717), .OUT(n4715) );
  NOR2 U2323 ( .A(n4719), .B(n4720), .OUT(n4718) );
  NOR2 U2324 ( .A(n4722), .B(n4723), .OUT(n4721) );
  NOR2 U2325 ( .A(n4725), .B(n4726), .OUT(n4724) );
  NOR2 U2326 ( .A(n4728), .B(n4729), .OUT(n4727) );
  NAND2 U2327 ( .A(n4731), .B(n4732), .OUT(n4730) );
  NOR2 U2328 ( .A(n4734), .B(n4735), .OUT(n4733) );
  NAND2 U2329 ( .A(n4737), .B(n4738), .OUT(n4736) );
  NAND2 U2330 ( .A(n4740), .B(n2028), .OUT(n4739) );
  NAND2 U2331 ( .A(n4742), .B(n2024), .OUT(n4741) );
  NAND2 U2332 ( .A(n4744), .B(n2020), .OUT(n4743) );
  NAND2 U2333 ( .A(n4746), .B(n2016), .OUT(n4745) );
  NAND2 U2334 ( .A(n4748), .B(n2012), .OUT(n4747) );
  NAND2 U2335 ( .A(n4750), .B(n2008), .OUT(n4749) );
  NAND2 U2336 ( .A(n4752), .B(n2004), .OUT(n4751) );
  NAND2 U2337 ( .A(n4754), .B(n2000), .OUT(n4753) );
  NAND2 U2338 ( .A(n4756), .B(n480), .OUT(n4755) );
  NAND2 U2339 ( .A(n4758), .B(n1996), .OUT(n4757) );
  NAND2 U2340 ( .A(n4760), .B(n1992), .OUT(n4759) );
  NAND2 U2341 ( .A(n4762), .B(n1988), .OUT(n4761) );
  NAND2 U2342 ( .A(n4764), .B(n1984), .OUT(n4763) );
  NAND2 U2343 ( .A(n4766), .B(n1980), .OUT(n4765) );
  NAND2 U2344 ( .A(n4768), .B(n1976), .OUT(n4767) );
  NAND2 U2345 ( .A(n4770), .B(n1972), .OUT(n4769) );
  NAND2 U2346 ( .A(n4772), .B(n1968), .OUT(n4771) );
  NAND2 U2347 ( .A(n4774), .B(n1964), .OUT(n4773) );
  NAND2 U2348 ( .A(n4776), .B(n1960), .OUT(n4775) );
  NAND2 U2349 ( .A(n4778), .B(n4779), .OUT(n4777) );
  NOR2 U2350 ( .A(n3802), .B(n2315), .OUT(n4780) );
  NAND2 U2351 ( .A(n2315), .B(n3802), .OUT(n4781) );
  NOR2 U2352 ( .A(n4780), .B(n4782), .OUT(\mult_49/A1[9] ) );
  NOR2 U2353 ( .A(n3806), .B(n2339), .OUT(n4783) );
  NAND2 U2354 ( .A(n2339), .B(n3806), .OUT(n4784) );
  NOR2 U2355 ( .A(n4783), .B(n4785), .OUT(\mult_49/A1[7] ) );
  NOR2 U2356 ( .A(n3810), .B(n2333), .OUT(n4786) );
  NAND2 U2357 ( .A(n2333), .B(n3810), .OUT(n4787) );
  NOR2 U2358 ( .A(n4786), .B(n4788), .OUT(\mult_49/A1[5] ) );
  NOR2 U2359 ( .A(n3814), .B(n2327), .OUT(n4789) );
  NAND2 U2360 ( .A(n2327), .B(n3814), .OUT(n4790) );
  NOR2 U2361 ( .A(n4789), .B(n4791), .OUT(\mult_49/A1[3] ) );
  NAND2 U2362 ( .A(n4498), .B(n4793), .OUT(n4792) );
  NAND2 U2363 ( .A(n4489), .B(n4795), .OUT(n4794) );
  NAND2 U2364 ( .A(n4492), .B(n4797), .OUT(n4796) );
  NAND2 U2365 ( .A(n4474), .B(n4799), .OUT(n4798) );
  NAND2 U2366 ( .A(n4495), .B(n4801), .OUT(n4800) );
  NAND2 U2367 ( .A(n4507), .B(n4803), .OUT(n4802) );
  NAND2 U2368 ( .A(n4465), .B(n4805), .OUT(n4804) );
  NAND2 U2369 ( .A(n4468), .B(n4807), .OUT(n4806) );
  NAND2 U2370 ( .A(n4450), .B(n4809), .OUT(n4808) );
  NAND2 U2371 ( .A(n4471), .B(n4811), .OUT(n4810) );
  NAND2 U2372 ( .A(n4483), .B(n4813), .OUT(n4812) );
  NAND2 U2373 ( .A(n4441), .B(n4815), .OUT(n4814) );
  NAND2 U2374 ( .A(n4444), .B(n4817), .OUT(n4816) );
  NAND2 U2375 ( .A(n4438), .B(n4819), .OUT(n4818) );
  NAND2 U2376 ( .A(\mult_49/ab[1][29] ), .B(\mult_49/ab[0][30] ), .OUT(n4820)
         );
  NAND2 U2377 ( .A(n4822), .B(n4823), .OUT(n4821) );
  NAND2 U2378 ( .A(n4435), .B(n4825), .OUT(n4824) );
  NAND2 U2379 ( .A(n4447), .B(n4827), .OUT(n4826) );
  NAND2 U2380 ( .A(n4459), .B(n4829), .OUT(n4828) );
  NAND2 U2381 ( .A(n4453), .B(n4831), .OUT(n4830) );
  NAND2 U2382 ( .A(n4456), .B(n4833), .OUT(n4832) );
  NAND2 U2383 ( .A(n4462), .B(n4835), .OUT(n4834) );
  NAND2 U2384 ( .A(n4477), .B(n4837), .OUT(n4836) );
  NAND2 U2385 ( .A(n4480), .B(n4839), .OUT(n4838) );
  NAND2 U2386 ( .A(n4486), .B(n4841), .OUT(n4840) );
  NAND2 U2387 ( .A(n4501), .B(n4843), .OUT(n4842) );
  NAND2 U2388 ( .A(n4504), .B(n4845), .OUT(n4844) );
  NAND2 U2389 ( .A(n4585), .B(n4847), .OUT(n4846) );
  NAND2 U2390 ( .A(n4738), .B(n4849), .OUT(n4848) );
  NAND2 U2391 ( .A(n4546), .B(n4851), .OUT(n4850) );
  NAND2 U2392 ( .A(n4733), .B(n4730), .OUT(n4852) );
  NOR2 U2393 ( .A(n4730), .B(n4733), .OUT(n4853) );
  NOR2 U2394 ( .A(n4854), .B(n4853), .OUT(\mult_49/A1[29] ) );
  NOR2 U2395 ( .A(n4739), .B(n3511), .OUT(n4855) );
  NAND2 U2396 ( .A(n3511), .B(n4739), .OUT(n4856) );
  NOR2 U2397 ( .A(n4855), .B(n4857), .OUT(\mult_49/A1[27] ) );
  NOR2 U2398 ( .A(n4743), .B(n3499), .OUT(n4858) );
  NAND2 U2399 ( .A(n3499), .B(n4743), .OUT(n4859) );
  NOR2 U2400 ( .A(n4858), .B(n4860), .OUT(\mult_49/A1[25] ) );
  NOR2 U2401 ( .A(n4747), .B(n3487), .OUT(n4861) );
  NAND2 U2402 ( .A(n3487), .B(n4747), .OUT(n4862) );
  NOR2 U2403 ( .A(n4861), .B(n4863), .OUT(\mult_49/A1[23] ) );
  NOR2 U2404 ( .A(n4751), .B(n3475), .OUT(n4864) );
  NAND2 U2405 ( .A(n3475), .B(n4751), .OUT(n4865) );
  NOR2 U2406 ( .A(n4864), .B(n4866), .OUT(\mult_49/A1[21] ) );
  NOR2 U2407 ( .A(n4755), .B(n2321), .OUT(n4867) );
  NOR2 U2408 ( .A(n4869), .B(n4870), .OUT(n4868) );
  NOR2 U2409 ( .A(n4867), .B(n4868), .OUT(\mult_49/A1[1] ) );
  NOR2 U2410 ( .A(n4757), .B(n3463), .OUT(n4871) );
  NAND2 U2411 ( .A(n3463), .B(n4757), .OUT(n4872) );
  NOR2 U2412 ( .A(n4871), .B(n4873), .OUT(\mult_49/A1[19] ) );
  NOR2 U2413 ( .A(n4761), .B(n3451), .OUT(n4874) );
  NAND2 U2414 ( .A(n3451), .B(n4761), .OUT(n4875) );
  NOR2 U2415 ( .A(n4874), .B(n4876), .OUT(\mult_49/A1[17] ) );
  NOR2 U2416 ( .A(n4765), .B(n3439), .OUT(n4877) );
  NAND2 U2417 ( .A(n3439), .B(n4765), .OUT(n4878) );
  NOR2 U2418 ( .A(n4877), .B(n4879), .OUT(\mult_49/A1[15] ) );
  NOR2 U2419 ( .A(n4769), .B(n3427), .OUT(n4880) );
  NAND2 U2420 ( .A(n3427), .B(n4769), .OUT(n4881) );
  NOR2 U2421 ( .A(n4880), .B(n4882), .OUT(\mult_49/A1[13] ) );
  NOR2 U2422 ( .A(n4773), .B(n3415), .OUT(n4883) );
  NAND2 U2423 ( .A(n3415), .B(n4773), .OUT(n4884) );
  NOR2 U2424 ( .A(n4883), .B(n4885), .OUT(\mult_49/A1[11] ) );
  NAND2 U2425 ( .A(n4887), .B(n4888), .OUT(n4886) );
  NOR2 U2426 ( .A(n3554), .B(n4886), .OUT(n4889) );
  NAND2 U2427 ( .A(n4886), .B(n3554), .OUT(n4890) );
  NOR2 U2428 ( .A(n4889), .B(n4891), .OUT(N99) );
  NAND2 U2429 ( .A(n4893), .B(n4894), .OUT(n4892) );
  NOR2 U2430 ( .A(n3557), .B(n4892), .OUT(n4895) );
  NAND2 U2431 ( .A(n4892), .B(n3557), .OUT(n4896) );
  NOR2 U2432 ( .A(n4895), .B(n4897), .OUT(N98) );
  NAND2 U2433 ( .A(n4899), .B(n4900), .OUT(n4898) );
  NOR2 U2434 ( .A(n3560), .B(n4898), .OUT(n4901) );
  NAND2 U2435 ( .A(n4898), .B(n3560), .OUT(n4902) );
  NOR2 U2436 ( .A(n4901), .B(n4903), .OUT(N97) );
  NAND2 U2437 ( .A(n4905), .B(n4906), .OUT(n4904) );
  NOR2 U2438 ( .A(n3563), .B(n4904), .OUT(n4907) );
  NAND2 U2439 ( .A(n4904), .B(n3563), .OUT(n4908) );
  NOR2 U2440 ( .A(n4907), .B(n4909), .OUT(N96) );
  NAND2 U2441 ( .A(n4911), .B(n4912), .OUT(n4910) );
  NOR2 U2442 ( .A(n3571), .B(n4910), .OUT(n4913) );
  NAND2 U2443 ( .A(n4910), .B(n3571), .OUT(n4914) );
  NOR2 U2444 ( .A(n4913), .B(n4915), .OUT(N95) );
  NAND2 U2445 ( .A(n4917), .B(n4918), .OUT(n4916) );
  NAND2 U2446 ( .A(n4920), .B(n4921), .OUT(n4919) );
  NOR2 U2447 ( .A(n4923), .B(n4919), .OUT(n4922) );
  NAND2 U2448 ( .A(n4919), .B(n4923), .OUT(n4924) );
  NOR2 U2449 ( .A(n4922), .B(n4925), .OUT(N124) );
  NAND2 U2450 ( .A(n4927), .B(n4928), .OUT(n4926) );
  NOR2 U2451 ( .A(n3568), .B(n4926), .OUT(n4929) );
  NAND2 U2452 ( .A(n4926), .B(n3568), .OUT(n4930) );
  NOR2 U2453 ( .A(n4929), .B(n4931), .OUT(N123) );
  NAND2 U2454 ( .A(n4933), .B(n4934), .OUT(n4932) );
  NOR2 U2455 ( .A(n3574), .B(n4932), .OUT(n4935) );
  NAND2 U2456 ( .A(n4932), .B(n3574), .OUT(n4936) );
  NOR2 U2457 ( .A(n4935), .B(n4937), .OUT(N122) );
  NAND2 U2458 ( .A(n4939), .B(n4940), .OUT(n4938) );
  NOR2 U2459 ( .A(n3577), .B(n4938), .OUT(n4941) );
  NAND2 U2460 ( .A(n4938), .B(n3577), .OUT(n4942) );
  NOR2 U2461 ( .A(n4941), .B(n4943), .OUT(N121) );
  NAND2 U2462 ( .A(n4945), .B(n4946), .OUT(n4944) );
  NOR2 U2463 ( .A(n3580), .B(n4944), .OUT(n4947) );
  NAND2 U2464 ( .A(n4944), .B(n3580), .OUT(n4948) );
  NOR2 U2465 ( .A(n4947), .B(n4949), .OUT(N120) );
  NAND2 U2466 ( .A(n4951), .B(n4952), .OUT(n4950) );
  NOR2 U2467 ( .A(n3583), .B(n4950), .OUT(n4953) );
  NAND2 U2468 ( .A(n4950), .B(n3583), .OUT(n4954) );
  NOR2 U2469 ( .A(n4953), .B(n4955), .OUT(N119) );
  NAND2 U2470 ( .A(n4957), .B(n4958), .OUT(n4956) );
  NOR2 U2471 ( .A(n3586), .B(n4956), .OUT(n4959) );
  NAND2 U2472 ( .A(n4956), .B(n3586), .OUT(n4960) );
  NOR2 U2473 ( .A(n4959), .B(n4961), .OUT(N118) );
  NAND2 U2474 ( .A(n4963), .B(n4964), .OUT(n4962) );
  NOR2 U2475 ( .A(n3589), .B(n4962), .OUT(n4965) );
  NAND2 U2476 ( .A(n4962), .B(n3589), .OUT(n4966) );
  NOR2 U2477 ( .A(n4965), .B(n4967), .OUT(N117) );
  NAND2 U2478 ( .A(n4969), .B(n4970), .OUT(n4968) );
  NOR2 U2479 ( .A(n3592), .B(n4968), .OUT(n4971) );
  NAND2 U2480 ( .A(n4968), .B(n3592), .OUT(n4972) );
  NOR2 U2481 ( .A(n4971), .B(n4973), .OUT(N116) );
  NAND2 U2482 ( .A(n4975), .B(n4976), .OUT(n4974) );
  NOR2 U2483 ( .A(n3595), .B(n4974), .OUT(n4977) );
  NAND2 U2484 ( .A(n4974), .B(n3595), .OUT(n4978) );
  NOR2 U2485 ( .A(n4977), .B(n4979), .OUT(N115) );
  NAND2 U2486 ( .A(n4981), .B(n4982), .OUT(n4980) );
  NOR2 U2487 ( .A(n3598), .B(n4980), .OUT(n4983) );
  NAND2 U2488 ( .A(n4980), .B(n3598), .OUT(n4984) );
  NOR2 U2489 ( .A(n4983), .B(n4985), .OUT(N114) );
  NAND2 U2490 ( .A(n4987), .B(n4988), .OUT(n4986) );
  NOR2 U2491 ( .A(n3601), .B(n4986), .OUT(n4989) );
  NAND2 U2492 ( .A(n4986), .B(n3601), .OUT(n4990) );
  NOR2 U2493 ( .A(n4989), .B(n4991), .OUT(N113) );
  NAND2 U2494 ( .A(n4993), .B(n4994), .OUT(n4992) );
  NOR2 U2495 ( .A(n3607), .B(n4992), .OUT(n4995) );
  NAND2 U2496 ( .A(n4992), .B(n3607), .OUT(n4996) );
  NOR2 U2497 ( .A(n4995), .B(n4997), .OUT(N112) );
  NAND2 U2498 ( .A(n4999), .B(n5000), .OUT(n4998) );
  NOR2 U2499 ( .A(n3610), .B(n4998), .OUT(n5001) );
  NAND2 U2500 ( .A(n4998), .B(n3610), .OUT(n5002) );
  NOR2 U2501 ( .A(n5001), .B(n5003), .OUT(N111) );
  NAND2 U2502 ( .A(n5005), .B(n5006), .OUT(n5004) );
  NOR2 U2503 ( .A(n3613), .B(n5004), .OUT(n5007) );
  NAND2 U2504 ( .A(n5004), .B(n3613), .OUT(n5008) );
  NOR2 U2505 ( .A(n5007), .B(n5009), .OUT(N110) );
  NAND2 U2506 ( .A(n5011), .B(n5012), .OUT(n5010) );
  NOR2 U2507 ( .A(n3616), .B(n5010), .OUT(n5013) );
  NAND2 U2508 ( .A(n5010), .B(n3616), .OUT(n5014) );
  NOR2 U2509 ( .A(n5013), .B(n5015), .OUT(N109) );
  NAND2 U2510 ( .A(n5017), .B(n5018), .OUT(n5016) );
  NOR2 U2511 ( .A(n3619), .B(n5016), .OUT(n5019) );
  NAND2 U2512 ( .A(n5016), .B(n3619), .OUT(n5020) );
  NOR2 U2513 ( .A(n5019), .B(n5021), .OUT(N108) );
  NAND2 U2514 ( .A(n5023), .B(n5024), .OUT(n5022) );
  NOR2 U2515 ( .A(n3622), .B(n5022), .OUT(n5025) );
  NAND2 U2516 ( .A(n5022), .B(n3622), .OUT(n5026) );
  NOR2 U2517 ( .A(n5025), .B(n5027), .OUT(N107) );
  NAND2 U2518 ( .A(n5029), .B(n5030), .OUT(n5028) );
  NOR2 U2519 ( .A(n3625), .B(n5028), .OUT(n5031) );
  NAND2 U2520 ( .A(n5028), .B(n3625), .OUT(n5032) );
  NOR2 U2521 ( .A(n5031), .B(n5033), .OUT(N106) );
  NAND2 U2522 ( .A(n5035), .B(n5036), .OUT(n5034) );
  NOR2 U2523 ( .A(n3628), .B(n5034), .OUT(n5037) );
  NAND2 U2524 ( .A(n5034), .B(n3628), .OUT(n5038) );
  NOR2 U2525 ( .A(n5037), .B(n5039), .OUT(N105) );
  NAND2 U2526 ( .A(n5041), .B(n5042), .OUT(n5040) );
  NOR2 U2527 ( .A(n3631), .B(n5040), .OUT(n5043) );
  NAND2 U2528 ( .A(n5040), .B(n3631), .OUT(n5044) );
  NOR2 U2529 ( .A(n5043), .B(n5045), .OUT(N104) );
  NAND2 U2530 ( .A(n5047), .B(n5048), .OUT(n5046) );
  NOR2 U2531 ( .A(n3634), .B(n5046), .OUT(n5049) );
  NAND2 U2532 ( .A(n5046), .B(n3634), .OUT(n5050) );
  NOR2 U2533 ( .A(n5049), .B(n5051), .OUT(N103) );
  NAND2 U2534 ( .A(n5053), .B(n5054), .OUT(n5052) );
  NOR2 U2535 ( .A(n3545), .B(n5052), .OUT(n5055) );
  NAND2 U2536 ( .A(n5052), .B(n3545), .OUT(n5056) );
  NOR2 U2537 ( .A(n5055), .B(n5057), .OUT(N102) );
  NAND2 U2538 ( .A(n5059), .B(n5060), .OUT(n5058) );
  NOR2 U2539 ( .A(n3548), .B(n5058), .OUT(n5061) );
  NAND2 U2540 ( .A(n5058), .B(n3548), .OUT(n5062) );
  NOR2 U2541 ( .A(n5061), .B(n5063), .OUT(N101) );
  NAND2 U2542 ( .A(n5065), .B(n5066), .OUT(n5064) );
  NOR2 U2543 ( .A(n3551), .B(n5064), .OUT(n5067) );
  NAND2 U2544 ( .A(n5064), .B(n3551), .OUT(n5068) );
  NOR2 U2545 ( .A(n5067), .B(n5069), .OUT(N100) );
  INV U2546 ( .IN(n1774), .OUT(n5070) );
  INV U2547 ( .IN(n1670), .OUT(n5071) );
  INV U2548 ( .IN(n1570), .OUT(n5072) );
  INV U2549 ( .IN(n1474), .OUT(n5073) );
  INV U2550 ( .IN(n1382), .OUT(n5074) );
  INV U2551 ( .IN(n1294), .OUT(n5075) );
  INV U2552 ( .IN(n1210), .OUT(n5076) );
  INV U2553 ( .IN(n1130), .OUT(n5077) );
  INV U2554 ( .IN(n1054), .OUT(n5078) );
  INV U2555 ( .IN(n982), .OUT(n5079) );
  INV U2556 ( .IN(n914), .OUT(n5080) );
  INV U2557 ( .IN(n850), .OUT(n5081) );
  INV U2558 ( .IN(n790), .OUT(n5082) );
  INV U2559 ( .IN(n734), .OUT(n5083) );
  INV U2560 ( .IN(n682), .OUT(n5084) );
  INV U2561 ( .IN(n634), .OUT(n5085) );
  INV U2562 ( .IN(n590), .OUT(n5086) );
  INV U2563 ( .IN(n550), .OUT(n5087) );
  INV U2564 ( .IN(n514), .OUT(n5088) );
  INV U2565 ( .IN(n291), .OUT(n5089) );
  INV U2566 ( .IN(n296), .OUT(n5090) );
  INV U2567 ( .IN(n304), .OUT(n5091) );
  INV U2568 ( .IN(n316), .OUT(n5092) );
  INV U2569 ( .IN(n332), .OUT(n5093) );
  INV U2570 ( .IN(n352), .OUT(n5094) );
  INV U2571 ( .IN(n376), .OUT(n5095) );
  INV U2572 ( .IN(n404), .OUT(n5096) );
  INV U2573 ( .IN(n436), .OUT(n5097) );
  INV U2574 ( .IN(n472), .OUT(n5098) );
  NAND2 U2575 ( .A(n5090), .B(n295), .OUT(n5099) );
  NAND2 U2576 ( .A(n2186), .B(n5099), .OUT(n302) );
  NAND2 U2577 ( .A(n296), .B(\mult_49/ab[2][8] ), .OUT(n301) );
  INV U2578 ( .IN(n300), .OUT(n5100) );
  NAND2 U2579 ( .A(n5091), .B(n303), .OUT(n5101) );
  NAND2 U2580 ( .A(n2192), .B(n5101), .OUT(n309) );
  NAND2 U2581 ( .A(n304), .B(\mult_49/ab[2][7] ), .OUT(n308) );
  INV U2582 ( .IN(n307), .OUT(n5102) );
  NAND2 U2583 ( .A(n5102), .B(n310), .OUT(n3770) );
  NAND2 U2584 ( .A(n2195), .B(n3770), .OUT(n314) );
  NAND2 U2585 ( .A(\mult_49/ab[3][7] ), .B(n307), .OUT(n313) );
  INV U2586 ( .IN(n312), .OUT(n5103) );
  NAND2 U2587 ( .A(n5092), .B(n315), .OUT(n5104) );
  NAND2 U2588 ( .A(n2201), .B(n5104), .OUT(n321) );
  NAND2 U2589 ( .A(n316), .B(\mult_49/ab[2][6] ), .OUT(n320) );
  INV U2590 ( .IN(n319), .OUT(n5105) );
  NAND2 U2591 ( .A(n5105), .B(n322), .OUT(n3755) );
  NAND2 U2592 ( .A(n2204), .B(n3755), .OUT(n325) );
  NAND2 U2593 ( .A(\mult_49/ab[3][6] ), .B(n319), .OUT(n324) );
  INV U2594 ( .IN(n323), .OUT(n5106) );
  NAND2 U2595 ( .A(n5106), .B(n326), .OUT(n3772) );
  NAND2 U2596 ( .A(n2207), .B(n3772), .OUT(n330) );
  NAND2 U2597 ( .A(\mult_49/ab[4][6] ), .B(n323), .OUT(n329) );
  INV U2598 ( .IN(n328), .OUT(n5107) );
  NAND2 U2599 ( .A(n5093), .B(n331), .OUT(n5108) );
  NAND2 U2600 ( .A(n2213), .B(n5108), .OUT(n337) );
  NAND2 U2601 ( .A(n332), .B(\mult_49/ab[2][5] ), .OUT(n336) );
  INV U2602 ( .IN(n335), .OUT(n5109) );
  NAND2 U2603 ( .A(n5109), .B(n338), .OUT(n3742) );
  NAND2 U2604 ( .A(n2216), .B(n3742), .OUT(n341) );
  NAND2 U2605 ( .A(\mult_49/ab[3][5] ), .B(n335), .OUT(n340) );
  INV U2606 ( .IN(n339), .OUT(n5110) );
  NAND2 U2607 ( .A(n5110), .B(n342), .OUT(n3757) );
  NAND2 U2608 ( .A(n2219), .B(n3757), .OUT(n345) );
  NAND2 U2609 ( .A(\mult_49/ab[4][5] ), .B(n339), .OUT(n344) );
  INV U2610 ( .IN(n343), .OUT(n5111) );
  NAND2 U2611 ( .A(n5111), .B(n346), .OUT(n3774) );
  NAND2 U2612 ( .A(n2222), .B(n3774), .OUT(n350) );
  NAND2 U2613 ( .A(\mult_49/ab[5][5] ), .B(n343), .OUT(n349) );
  INV U2614 ( .IN(n348), .OUT(n5112) );
  NAND2 U2615 ( .A(n5094), .B(n351), .OUT(n5113) );
  NAND2 U2616 ( .A(n2228), .B(n5113), .OUT(n357) );
  NAND2 U2617 ( .A(n352), .B(\mult_49/ab[2][4] ), .OUT(n356) );
  INV U2618 ( .IN(n355), .OUT(n5114) );
  NAND2 U2619 ( .A(n5114), .B(n358), .OUT(n3731) );
  NAND2 U2620 ( .A(n2231), .B(n3731), .OUT(n361) );
  NAND2 U2621 ( .A(\mult_49/ab[3][4] ), .B(n355), .OUT(n360) );
  INV U2622 ( .IN(n359), .OUT(n5115) );
  NAND2 U2623 ( .A(n5115), .B(n362), .OUT(n3744) );
  NAND2 U2624 ( .A(n2234), .B(n3744), .OUT(n365) );
  NAND2 U2625 ( .A(\mult_49/ab[4][4] ), .B(n359), .OUT(n364) );
  INV U2626 ( .IN(n363), .OUT(n5116) );
  NAND2 U2627 ( .A(n5116), .B(n366), .OUT(n3759) );
  NAND2 U2628 ( .A(n2237), .B(n3759), .OUT(n369) );
  NAND2 U2629 ( .A(\mult_49/ab[5][4] ), .B(n363), .OUT(n368) );
  INV U2630 ( .IN(n367), .OUT(n5117) );
  NAND2 U2631 ( .A(n5117), .B(n370), .OUT(n3776) );
  NAND2 U2632 ( .A(n2240), .B(n3776), .OUT(n374) );
  NAND2 U2633 ( .A(\mult_49/ab[6][4] ), .B(n367), .OUT(n373) );
  INV U2634 ( .IN(n372), .OUT(n5118) );
  NAND2 U2635 ( .A(n5095), .B(n375), .OUT(n5119) );
  NAND2 U2636 ( .A(n2246), .B(n5119), .OUT(n381) );
  NAND2 U2637 ( .A(n376), .B(\mult_49/ab[2][3] ), .OUT(n380) );
  INV U2638 ( .IN(n379), .OUT(n5120) );
  NAND2 U2639 ( .A(n5120), .B(n382), .OUT(n3722) );
  NAND2 U2640 ( .A(n2249), .B(n3722), .OUT(n385) );
  NAND2 U2641 ( .A(\mult_49/ab[3][3] ), .B(n379), .OUT(n384) );
  INV U2642 ( .IN(n383), .OUT(n5121) );
  NAND2 U2643 ( .A(n5121), .B(n386), .OUT(n3733) );
  NAND2 U2644 ( .A(n2252), .B(n3733), .OUT(n389) );
  NAND2 U2645 ( .A(\mult_49/ab[4][3] ), .B(n383), .OUT(n388) );
  INV U2646 ( .IN(n387), .OUT(n5122) );
  NAND2 U2647 ( .A(n5122), .B(n390), .OUT(n3746) );
  NAND2 U2648 ( .A(n2255), .B(n3746), .OUT(n393) );
  NAND2 U2649 ( .A(\mult_49/ab[5][3] ), .B(n387), .OUT(n392) );
  INV U2650 ( .IN(n391), .OUT(n5123) );
  NAND2 U2651 ( .A(n5123), .B(n394), .OUT(n3761) );
  NAND2 U2652 ( .A(n2258), .B(n3761), .OUT(n397) );
  NAND2 U2653 ( .A(\mult_49/ab[6][3] ), .B(n391), .OUT(n396) );
  INV U2654 ( .IN(n395), .OUT(n5124) );
  NAND2 U2655 ( .A(n5124), .B(n398), .OUT(n3778) );
  NAND2 U2656 ( .A(n2261), .B(n3778), .OUT(n402) );
  NAND2 U2657 ( .A(\mult_49/ab[7][3] ), .B(n395), .OUT(n401) );
  INV U2658 ( .IN(n400), .OUT(n5125) );
  NAND2 U2659 ( .A(n5096), .B(n403), .OUT(n5126) );
  NAND2 U2660 ( .A(n2267), .B(n5126), .OUT(n409) );
  NAND2 U2661 ( .A(n404), .B(\mult_49/ab[2][2] ), .OUT(n408) );
  INV U2662 ( .IN(n407), .OUT(n5127) );
  NAND2 U2663 ( .A(n5127), .B(n410), .OUT(n3715) );
  NAND2 U2664 ( .A(n2270), .B(n3715), .OUT(n413) );
  NAND2 U2665 ( .A(\mult_49/ab[3][2] ), .B(n407), .OUT(n412) );
  INV U2666 ( .IN(n411), .OUT(n5128) );
  NAND2 U2667 ( .A(n5128), .B(n414), .OUT(n3724) );
  NAND2 U2668 ( .A(n2273), .B(n3724), .OUT(n417) );
  NAND2 U2669 ( .A(\mult_49/ab[4][2] ), .B(n411), .OUT(n416) );
  INV U2670 ( .IN(n415), .OUT(n5129) );
  NAND2 U2671 ( .A(n5129), .B(n418), .OUT(n3735) );
  NAND2 U2672 ( .A(n2276), .B(n3735), .OUT(n421) );
  NAND2 U2673 ( .A(\mult_49/ab[5][2] ), .B(n415), .OUT(n420) );
  INV U2674 ( .IN(n419), .OUT(n5130) );
  NAND2 U2675 ( .A(n5130), .B(n422), .OUT(n3748) );
  NAND2 U2676 ( .A(n2279), .B(n3748), .OUT(n425) );
  NAND2 U2677 ( .A(\mult_49/ab[6][2] ), .B(n419), .OUT(n424) );
  INV U2678 ( .IN(n423), .OUT(n5131) );
  NAND2 U2679 ( .A(n5131), .B(n426), .OUT(n3763) );
  NAND2 U2680 ( .A(n2282), .B(n3763), .OUT(n429) );
  NAND2 U2681 ( .A(\mult_49/ab[7][2] ), .B(n423), .OUT(n428) );
  INV U2682 ( .IN(n427), .OUT(n5132) );
  NAND2 U2683 ( .A(n5132), .B(n430), .OUT(n3780) );
  NAND2 U2684 ( .A(n2285), .B(n3780), .OUT(n434) );
  NAND2 U2685 ( .A(\mult_49/ab[8][2] ), .B(n427), .OUT(n433) );
  INV U2686 ( .IN(n432), .OUT(n5133) );
  NAND2 U2687 ( .A(n5097), .B(n435), .OUT(n5134) );
  NAND2 U2688 ( .A(n2291), .B(n5134), .OUT(n441) );
  NAND2 U2689 ( .A(n436), .B(\mult_49/ab[2][1] ), .OUT(n440) );
  INV U2690 ( .IN(n439), .OUT(n5135) );
  NAND2 U2691 ( .A(n5135), .B(n442), .OUT(n3710) );
  NAND2 U2692 ( .A(n2294), .B(n3710), .OUT(n445) );
  NAND2 U2693 ( .A(\mult_49/ab[3][1] ), .B(n439), .OUT(n444) );
  INV U2694 ( .IN(n443), .OUT(n5136) );
  NAND2 U2695 ( .A(n5136), .B(n446), .OUT(n3717) );
  NAND2 U2696 ( .A(n2297), .B(n3717), .OUT(n449) );
  NAND2 U2697 ( .A(\mult_49/ab[4][1] ), .B(n443), .OUT(n448) );
  INV U2698 ( .IN(n447), .OUT(n5137) );
  NAND2 U2699 ( .A(n5137), .B(n450), .OUT(n3726) );
  NAND2 U2700 ( .A(n2300), .B(n3726), .OUT(n453) );
  NAND2 U2701 ( .A(\mult_49/ab[5][1] ), .B(n447), .OUT(n452) );
  INV U2702 ( .IN(n451), .OUT(n5138) );
  NAND2 U2703 ( .A(n5138), .B(n454), .OUT(n3737) );
  NAND2 U2704 ( .A(n2303), .B(n3737), .OUT(n457) );
  NAND2 U2705 ( .A(\mult_49/ab[6][1] ), .B(n451), .OUT(n456) );
  INV U2706 ( .IN(n455), .OUT(n5139) );
  NAND2 U2707 ( .A(n5139), .B(n458), .OUT(n3750) );
  NAND2 U2708 ( .A(n2306), .B(n3750), .OUT(n461) );
  NAND2 U2709 ( .A(\mult_49/ab[7][1] ), .B(n455), .OUT(n460) );
  INV U2710 ( .IN(n459), .OUT(n5140) );
  NAND2 U2711 ( .A(n5140), .B(n462), .OUT(n3765) );
  NAND2 U2712 ( .A(n2309), .B(n3765), .OUT(n465) );
  NAND2 U2713 ( .A(\mult_49/ab[8][1] ), .B(n459), .OUT(n464) );
  INV U2714 ( .IN(n463), .OUT(n5141) );
  NAND2 U2715 ( .A(n5141), .B(n466), .OUT(n3782) );
  NAND2 U2716 ( .A(n2312), .B(n3782), .OUT(n470) );
  NAND2 U2717 ( .A(\mult_49/ab[9][1] ), .B(n463), .OUT(n469) );
  INV U2718 ( .IN(n468), .OUT(n5142) );
  NAND2 U2719 ( .A(n5098), .B(n471), .OUT(n5143) );
  NAND2 U2720 ( .A(n2318), .B(n5143), .OUT(n477) );
  NAND2 U2721 ( .A(n472), .B(\mult_49/ab[2][0] ), .OUT(n476) );
  INV U2722 ( .IN(n475), .OUT(n5144) );
  NAND2 U2723 ( .A(n4869), .B(n4756), .OUT(n481) );
  INV U2724 ( .IN(n479), .OUT(n5145) );
  NAND2 U2725 ( .A(n2324), .B(n3817), .OUT(n485) );
  INV U2726 ( .IN(n483), .OUT(n5146) );
  NAND2 U2727 ( .A(n5147), .B(n3815), .OUT(n489) );
  INV U2728 ( .IN(n487), .OUT(n5148) );
  NAND2 U2729 ( .A(n2330), .B(n3813), .OUT(n493) );
  INV U2730 ( .IN(n491), .OUT(n5149) );
  NAND2 U2731 ( .A(n5150), .B(n3811), .OUT(n497) );
  INV U2732 ( .IN(n495), .OUT(n5151) );
  NAND2 U2733 ( .A(n2336), .B(n3809), .OUT(n501) );
  INV U2734 ( .IN(n499), .OUT(n5152) );
  NAND2 U2735 ( .A(n5153), .B(n3807), .OUT(n505) );
  INV U2736 ( .IN(n503), .OUT(n5154) );
  NAND2 U2737 ( .A(n2342), .B(n3805), .OUT(n510) );
  INV U2738 ( .IN(n508), .OUT(n5155) );
  NAND2 U2739 ( .A(n5070), .B(n1777), .OUT(n5156) );
  NAND2 U2740 ( .A(n5157), .B(n5156), .OUT(n4823) );
  NAND2 U2741 ( .A(\mult_49/ab[2][28] ), .B(n1774), .OUT(n4822) );
  NAND2 U2742 ( .A(n5071), .B(n1673), .OUT(n5158) );
  NAND2 U2743 ( .A(n3220), .B(n5158), .OUT(n1781) );
  NAND2 U2744 ( .A(\mult_49/ab[2][27] ), .B(n1670), .OUT(n1780) );
  INV U2745 ( .IN(n1779), .OUT(n5159) );
  NAND2 U2746 ( .A(n5159), .B(n1778), .OUT(n4434) );
  NAND2 U2747 ( .A(n3301), .B(n4434), .OUT(n4825) );
  NAND2 U2748 ( .A(\mult_49/ab[3][27] ), .B(n1779), .OUT(n4435) );
  NAND2 U2749 ( .A(n5072), .B(n1573), .OUT(n5160) );
  NAND2 U2750 ( .A(n3145), .B(n5160), .OUT(n1677) );
  NAND2 U2751 ( .A(\mult_49/ab[2][26] ), .B(n1570), .OUT(n1676) );
  INV U2752 ( .IN(n1675), .OUT(n5161) );
  NAND2 U2753 ( .A(n5161), .B(n1674), .OUT(n4383) );
  NAND2 U2754 ( .A(n3223), .B(n4383), .OUT(n1785) );
  NAND2 U2755 ( .A(\mult_49/ab[3][26] ), .B(n1675), .OUT(n1784) );
  INV U2756 ( .IN(n1783), .OUT(n5162) );
  NAND2 U2757 ( .A(n5162), .B(n1782), .OUT(n4437) );
  NAND2 U2758 ( .A(n3304), .B(n4437), .OUT(n4819) );
  NAND2 U2759 ( .A(\mult_49/ab[4][26] ), .B(n1783), .OUT(n4438) );
  NAND2 U2760 ( .A(n5073), .B(n1477), .OUT(n5163) );
  NAND2 U2761 ( .A(n3073), .B(n5163), .OUT(n1577) );
  NAND2 U2762 ( .A(\mult_49/ab[2][25] ), .B(n1474), .OUT(n1576) );
  INV U2763 ( .IN(n1575), .OUT(n5164) );
  NAND2 U2764 ( .A(n5164), .B(n1574), .OUT(n4334) );
  NAND2 U2765 ( .A(n3148), .B(n4334), .OUT(n1681) );
  NAND2 U2766 ( .A(\mult_49/ab[3][25] ), .B(n1575), .OUT(n1680) );
  INV U2767 ( .IN(n1679), .OUT(n5165) );
  NAND2 U2768 ( .A(n5165), .B(n1678), .OUT(n4385) );
  NAND2 U2769 ( .A(n3226), .B(n4385), .OUT(n1789) );
  NAND2 U2770 ( .A(\mult_49/ab[4][25] ), .B(n1679), .OUT(n1788) );
  INV U2771 ( .IN(n1787), .OUT(n5166) );
  NAND2 U2772 ( .A(n5166), .B(n1786), .OUT(n4440) );
  NAND2 U2773 ( .A(n3307), .B(n4440), .OUT(n4815) );
  NAND2 U2774 ( .A(\mult_49/ab[5][25] ), .B(n1787), .OUT(n4441) );
  NAND2 U2775 ( .A(n5074), .B(n1385), .OUT(n5167) );
  NAND2 U2776 ( .A(n3004), .B(n5167), .OUT(n1481) );
  NAND2 U2777 ( .A(\mult_49/ab[2][24] ), .B(n1382), .OUT(n1480) );
  INV U2778 ( .IN(n1479), .OUT(n5168) );
  NAND2 U2779 ( .A(n5168), .B(n1478), .OUT(n4287) );
  NAND2 U2780 ( .A(n3076), .B(n4287), .OUT(n1581) );
  NAND2 U2781 ( .A(\mult_49/ab[3][24] ), .B(n1479), .OUT(n1580) );
  INV U2782 ( .IN(n1579), .OUT(n5169) );
  NAND2 U2783 ( .A(n5169), .B(n1578), .OUT(n4336) );
  NAND2 U2784 ( .A(n3151), .B(n4336), .OUT(n1685) );
  NAND2 U2785 ( .A(\mult_49/ab[4][24] ), .B(n1579), .OUT(n1684) );
  INV U2786 ( .IN(n1683), .OUT(n5170) );
  NAND2 U2787 ( .A(n5170), .B(n1682), .OUT(n4387) );
  NAND2 U2788 ( .A(n3229), .B(n4387), .OUT(n1793) );
  NAND2 U2789 ( .A(\mult_49/ab[5][24] ), .B(n1683), .OUT(n1792) );
  INV U2790 ( .IN(n1791), .OUT(n5171) );
  NAND2 U2791 ( .A(n5171), .B(n1790), .OUT(n4443) );
  NAND2 U2792 ( .A(n3310), .B(n4443), .OUT(n4817) );
  NAND2 U2793 ( .A(\mult_49/ab[6][24] ), .B(n1791), .OUT(n4444) );
  NAND2 U2794 ( .A(n5075), .B(n1297), .OUT(n5172) );
  NAND2 U2795 ( .A(n2938), .B(n5172), .OUT(n1389) );
  NAND2 U2796 ( .A(\mult_49/ab[2][23] ), .B(n1294), .OUT(n1388) );
  INV U2797 ( .IN(n1387), .OUT(n5173) );
  NAND2 U2798 ( .A(n5173), .B(n1386), .OUT(n4242) );
  NAND2 U2799 ( .A(n3007), .B(n4242), .OUT(n1485) );
  NAND2 U2800 ( .A(\mult_49/ab[3][23] ), .B(n1387), .OUT(n1484) );
  INV U2801 ( .IN(n1483), .OUT(n5174) );
  NAND2 U2802 ( .A(n5174), .B(n1482), .OUT(n4289) );
  NAND2 U2803 ( .A(n3079), .B(n4289), .OUT(n1585) );
  NAND2 U2804 ( .A(\mult_49/ab[4][23] ), .B(n1483), .OUT(n1584) );
  INV U2805 ( .IN(n1583), .OUT(n5175) );
  NAND2 U2806 ( .A(n5175), .B(n1582), .OUT(n4338) );
  NAND2 U2807 ( .A(n3154), .B(n4338), .OUT(n1689) );
  NAND2 U2808 ( .A(\mult_49/ab[5][23] ), .B(n1583), .OUT(n1688) );
  INV U2809 ( .IN(n1687), .OUT(n5176) );
  NAND2 U2810 ( .A(n5176), .B(n1686), .OUT(n4389) );
  NAND2 U2811 ( .A(n3232), .B(n4389), .OUT(n1797) );
  NAND2 U2812 ( .A(\mult_49/ab[6][23] ), .B(n1687), .OUT(n1796) );
  INV U2813 ( .IN(n1795), .OUT(n5177) );
  NAND2 U2814 ( .A(n5177), .B(n1794), .OUT(n4446) );
  NAND2 U2815 ( .A(n3313), .B(n4446), .OUT(n4827) );
  NAND2 U2816 ( .A(\mult_49/ab[7][23] ), .B(n1795), .OUT(n4447) );
  NAND2 U2817 ( .A(n5076), .B(n1213), .OUT(n5178) );
  NAND2 U2818 ( .A(n2875), .B(n5178), .OUT(n1301) );
  NAND2 U2819 ( .A(\mult_49/ab[2][22] ), .B(n1210), .OUT(n1300) );
  INV U2820 ( .IN(n1299), .OUT(n5179) );
  NAND2 U2821 ( .A(n5179), .B(n1298), .OUT(n4199) );
  NAND2 U2822 ( .A(n2941), .B(n4199), .OUT(n1393) );
  NAND2 U2823 ( .A(\mult_49/ab[3][22] ), .B(n1299), .OUT(n1392) );
  INV U2824 ( .IN(n1391), .OUT(n5180) );
  NAND2 U2825 ( .A(n5180), .B(n1390), .OUT(n4244) );
  NAND2 U2826 ( .A(n3010), .B(n4244), .OUT(n1489) );
  NAND2 U2827 ( .A(\mult_49/ab[4][22] ), .B(n1391), .OUT(n1488) );
  INV U2828 ( .IN(n1487), .OUT(n5181) );
  NAND2 U2829 ( .A(n5181), .B(n1486), .OUT(n4291) );
  NAND2 U2830 ( .A(n3082), .B(n4291), .OUT(n1589) );
  NAND2 U2831 ( .A(\mult_49/ab[5][22] ), .B(n1487), .OUT(n1588) );
  INV U2832 ( .IN(n1587), .OUT(n5182) );
  NAND2 U2833 ( .A(n5182), .B(n1586), .OUT(n4340) );
  NAND2 U2834 ( .A(n3157), .B(n4340), .OUT(n1693) );
  NAND2 U2835 ( .A(\mult_49/ab[6][22] ), .B(n1587), .OUT(n1692) );
  INV U2836 ( .IN(n1691), .OUT(n5183) );
  NAND2 U2837 ( .A(n5183), .B(n1690), .OUT(n4391) );
  NAND2 U2838 ( .A(n3235), .B(n4391), .OUT(n1801) );
  NAND2 U2839 ( .A(\mult_49/ab[7][22] ), .B(n1691), .OUT(n1800) );
  INV U2840 ( .IN(n1799), .OUT(n5184) );
  NAND2 U2841 ( .A(n5184), .B(n1798), .OUT(n4449) );
  NAND2 U2842 ( .A(n3316), .B(n4449), .OUT(n4809) );
  NAND2 U2843 ( .A(\mult_49/ab[8][22] ), .B(n1799), .OUT(n4450) );
  NAND2 U2844 ( .A(n5077), .B(n1133), .OUT(n5185) );
  NAND2 U2845 ( .A(n2815), .B(n5185), .OUT(n1217) );
  NAND2 U2846 ( .A(\mult_49/ab[2][21] ), .B(n1130), .OUT(n1216) );
  INV U2847 ( .IN(n1215), .OUT(n5186) );
  NAND2 U2848 ( .A(n5186), .B(n1214), .OUT(n4158) );
  NAND2 U2849 ( .A(n2878), .B(n4158), .OUT(n1305) );
  NAND2 U2850 ( .A(\mult_49/ab[3][21] ), .B(n1215), .OUT(n1304) );
  INV U2851 ( .IN(n1303), .OUT(n5187) );
  NAND2 U2852 ( .A(n5187), .B(n1302), .OUT(n4201) );
  NAND2 U2853 ( .A(n2944), .B(n4201), .OUT(n1397) );
  NAND2 U2854 ( .A(\mult_49/ab[4][21] ), .B(n1303), .OUT(n1396) );
  INV U2855 ( .IN(n1395), .OUT(n5188) );
  NAND2 U2856 ( .A(n5188), .B(n1394), .OUT(n4246) );
  NAND2 U2857 ( .A(n3013), .B(n4246), .OUT(n1493) );
  NAND2 U2858 ( .A(\mult_49/ab[5][21] ), .B(n1395), .OUT(n1492) );
  INV U2859 ( .IN(n1491), .OUT(n5189) );
  NAND2 U2860 ( .A(n5189), .B(n1490), .OUT(n4293) );
  NAND2 U2861 ( .A(n3085), .B(n4293), .OUT(n1593) );
  NAND2 U2862 ( .A(\mult_49/ab[6][21] ), .B(n1491), .OUT(n1592) );
  INV U2863 ( .IN(n1591), .OUT(n5190) );
  NAND2 U2864 ( .A(n5190), .B(n1590), .OUT(n4342) );
  NAND2 U2865 ( .A(n3160), .B(n4342), .OUT(n1697) );
  NAND2 U2866 ( .A(\mult_49/ab[7][21] ), .B(n1591), .OUT(n1696) );
  INV U2867 ( .IN(n1695), .OUT(n5191) );
  NAND2 U2868 ( .A(n5191), .B(n1694), .OUT(n4393) );
  NAND2 U2869 ( .A(n3238), .B(n4393), .OUT(n1805) );
  NAND2 U2870 ( .A(\mult_49/ab[8][21] ), .B(n1695), .OUT(n1804) );
  INV U2871 ( .IN(n1803), .OUT(n5192) );
  NAND2 U2872 ( .A(n5192), .B(n1802), .OUT(n4452) );
  NAND2 U2873 ( .A(n3319), .B(n4452), .OUT(n4831) );
  NAND2 U2874 ( .A(\mult_49/ab[9][21] ), .B(n1803), .OUT(n4453) );
  NAND2 U2875 ( .A(n5078), .B(n1057), .OUT(n5193) );
  NAND2 U2876 ( .A(n2758), .B(n5193), .OUT(n1137) );
  NAND2 U2877 ( .A(\mult_49/ab[2][20] ), .B(n1054), .OUT(n1136) );
  INV U2878 ( .IN(n1135), .OUT(n5194) );
  NAND2 U2879 ( .A(n5194), .B(n1134), .OUT(n4119) );
  NAND2 U2880 ( .A(n2818), .B(n4119), .OUT(n1221) );
  NAND2 U2881 ( .A(\mult_49/ab[3][20] ), .B(n1135), .OUT(n1220) );
  INV U2882 ( .IN(n1219), .OUT(n5195) );
  NAND2 U2883 ( .A(n5195), .B(n1218), .OUT(n4160) );
  NAND2 U2884 ( .A(n2881), .B(n4160), .OUT(n1309) );
  NAND2 U2885 ( .A(\mult_49/ab[4][20] ), .B(n1219), .OUT(n1308) );
  INV U2886 ( .IN(n1307), .OUT(n5196) );
  NAND2 U2887 ( .A(n5196), .B(n1306), .OUT(n4203) );
  NAND2 U2888 ( .A(n2947), .B(n4203), .OUT(n1401) );
  NAND2 U2889 ( .A(\mult_49/ab[5][20] ), .B(n1307), .OUT(n1400) );
  INV U2890 ( .IN(n1399), .OUT(n5197) );
  NAND2 U2891 ( .A(n5197), .B(n1398), .OUT(n4248) );
  NAND2 U2892 ( .A(n3016), .B(n4248), .OUT(n1497) );
  NAND2 U2893 ( .A(\mult_49/ab[6][20] ), .B(n1399), .OUT(n1496) );
  INV U2894 ( .IN(n1495), .OUT(n5198) );
  NAND2 U2895 ( .A(n5198), .B(n1494), .OUT(n4295) );
  NAND2 U2896 ( .A(n3088), .B(n4295), .OUT(n1597) );
  NAND2 U2897 ( .A(\mult_49/ab[7][20] ), .B(n1495), .OUT(n1596) );
  INV U2898 ( .IN(n1595), .OUT(n5199) );
  NAND2 U2899 ( .A(n5199), .B(n1594), .OUT(n4344) );
  NAND2 U2900 ( .A(n3163), .B(n4344), .OUT(n1701) );
  NAND2 U2901 ( .A(\mult_49/ab[8][20] ), .B(n1595), .OUT(n1700) );
  INV U2902 ( .IN(n1699), .OUT(n5200) );
  NAND2 U2903 ( .A(n5200), .B(n1698), .OUT(n4395) );
  NAND2 U2904 ( .A(n3241), .B(n4395), .OUT(n1809) );
  NAND2 U2905 ( .A(\mult_49/ab[9][20] ), .B(n1699), .OUT(n1808) );
  INV U2906 ( .IN(n1807), .OUT(n5201) );
  NAND2 U2907 ( .A(n5201), .B(n1806), .OUT(n4455) );
  NAND2 U2908 ( .A(n3322), .B(n4455), .OUT(n4833) );
  NAND2 U2909 ( .A(\mult_49/ab[10][20] ), .B(n1807), .OUT(n4456) );
  NAND2 U2910 ( .A(n5079), .B(n985), .OUT(n5202) );
  NAND2 U2911 ( .A(n2704), .B(n5202), .OUT(n1061) );
  NAND2 U2912 ( .A(\mult_49/ab[2][19] ), .B(n982), .OUT(n1060) );
  INV U2913 ( .IN(n1059), .OUT(n5203) );
  NAND2 U2914 ( .A(n5203), .B(n1058), .OUT(n4082) );
  NAND2 U2915 ( .A(n2761), .B(n4082), .OUT(n1141) );
  NAND2 U2916 ( .A(\mult_49/ab[3][19] ), .B(n1059), .OUT(n1140) );
  INV U2917 ( .IN(n1139), .OUT(n5204) );
  NAND2 U2918 ( .A(n5204), .B(n1138), .OUT(n4121) );
  NAND2 U2919 ( .A(n2821), .B(n4121), .OUT(n1225) );
  NAND2 U2920 ( .A(\mult_49/ab[4][19] ), .B(n1139), .OUT(n1224) );
  INV U2921 ( .IN(n1223), .OUT(n5205) );
  NAND2 U2922 ( .A(n5205), .B(n1222), .OUT(n4162) );
  NAND2 U2923 ( .A(n2884), .B(n4162), .OUT(n1313) );
  NAND2 U2924 ( .A(\mult_49/ab[5][19] ), .B(n1223), .OUT(n1312) );
  INV U2925 ( .IN(n1311), .OUT(n5206) );
  NAND2 U2926 ( .A(n5206), .B(n1310), .OUT(n4205) );
  NAND2 U2927 ( .A(n2950), .B(n4205), .OUT(n1405) );
  NAND2 U2928 ( .A(\mult_49/ab[6][19] ), .B(n1311), .OUT(n1404) );
  INV U2929 ( .IN(n1403), .OUT(n5207) );
  NAND2 U2930 ( .A(n5207), .B(n1402), .OUT(n4250) );
  NAND2 U2931 ( .A(n3019), .B(n4250), .OUT(n1501) );
  NAND2 U2932 ( .A(\mult_49/ab[7][19] ), .B(n1403), .OUT(n1500) );
  INV U2933 ( .IN(n1499), .OUT(n5208) );
  NAND2 U2934 ( .A(n5208), .B(n1498), .OUT(n4297) );
  NAND2 U2935 ( .A(n3091), .B(n4297), .OUT(n1601) );
  NAND2 U2936 ( .A(\mult_49/ab[8][19] ), .B(n1499), .OUT(n1600) );
  INV U2937 ( .IN(n1599), .OUT(n5209) );
  NAND2 U2938 ( .A(n5209), .B(n1598), .OUT(n4346) );
  NAND2 U2939 ( .A(n3166), .B(n4346), .OUT(n1705) );
  NAND2 U2940 ( .A(\mult_49/ab[9][19] ), .B(n1599), .OUT(n1704) );
  INV U2941 ( .IN(n1703), .OUT(n5210) );
  NAND2 U2942 ( .A(n5210), .B(n1702), .OUT(n4397) );
  NAND2 U2943 ( .A(n3244), .B(n4397), .OUT(n1813) );
  NAND2 U2944 ( .A(\mult_49/ab[10][19] ), .B(n1703), .OUT(n1812) );
  INV U2945 ( .IN(n1811), .OUT(n5211) );
  NAND2 U2946 ( .A(n5211), .B(n1810), .OUT(n4458) );
  NAND2 U2947 ( .A(n3325), .B(n4458), .OUT(n4829) );
  NAND2 U2948 ( .A(\mult_49/ab[11][19] ), .B(n1811), .OUT(n4459) );
  NAND2 U2949 ( .A(n5080), .B(n917), .OUT(n5212) );
  NAND2 U2950 ( .A(n2653), .B(n5212), .OUT(n989) );
  NAND2 U2951 ( .A(\mult_49/ab[2][18] ), .B(n914), .OUT(n988) );
  INV U2952 ( .IN(n987), .OUT(n5213) );
  NAND2 U2953 ( .A(n5213), .B(n986), .OUT(n4047) );
  NAND2 U2954 ( .A(n2707), .B(n4047), .OUT(n1065) );
  NAND2 U2955 ( .A(\mult_49/ab[3][18] ), .B(n987), .OUT(n1064) );
  INV U2956 ( .IN(n1063), .OUT(n5214) );
  NAND2 U2957 ( .A(n5214), .B(n1062), .OUT(n4084) );
  NAND2 U2958 ( .A(n2764), .B(n4084), .OUT(n1145) );
  NAND2 U2959 ( .A(\mult_49/ab[4][18] ), .B(n1063), .OUT(n1144) );
  INV U2960 ( .IN(n1143), .OUT(n5215) );
  NAND2 U2961 ( .A(n5215), .B(n1142), .OUT(n4123) );
  NAND2 U2962 ( .A(n2824), .B(n4123), .OUT(n1229) );
  NAND2 U2963 ( .A(\mult_49/ab[5][18] ), .B(n1143), .OUT(n1228) );
  INV U2964 ( .IN(n1227), .OUT(n5216) );
  NAND2 U2965 ( .A(n5216), .B(n1226), .OUT(n4164) );
  NAND2 U2966 ( .A(n2887), .B(n4164), .OUT(n1317) );
  NAND2 U2967 ( .A(\mult_49/ab[6][18] ), .B(n1227), .OUT(n1316) );
  INV U2968 ( .IN(n1315), .OUT(n5217) );
  NAND2 U2969 ( .A(n5217), .B(n1314), .OUT(n4207) );
  NAND2 U2970 ( .A(n2953), .B(n4207), .OUT(n1409) );
  NAND2 U2971 ( .A(\mult_49/ab[7][18] ), .B(n1315), .OUT(n1408) );
  INV U2972 ( .IN(n1407), .OUT(n5218) );
  NAND2 U2973 ( .A(n5218), .B(n1406), .OUT(n4252) );
  NAND2 U2974 ( .A(n3022), .B(n4252), .OUT(n1505) );
  NAND2 U2975 ( .A(\mult_49/ab[8][18] ), .B(n1407), .OUT(n1504) );
  INV U2976 ( .IN(n1503), .OUT(n5219) );
  NAND2 U2977 ( .A(n5219), .B(n1502), .OUT(n4299) );
  NAND2 U2978 ( .A(n3094), .B(n4299), .OUT(n1605) );
  NAND2 U2979 ( .A(\mult_49/ab[9][18] ), .B(n1503), .OUT(n1604) );
  INV U2980 ( .IN(n1603), .OUT(n5220) );
  NAND2 U2981 ( .A(n5220), .B(n1602), .OUT(n4348) );
  NAND2 U2982 ( .A(n3169), .B(n4348), .OUT(n1709) );
  NAND2 U2983 ( .A(\mult_49/ab[10][18] ), .B(n1603), .OUT(n1708) );
  INV U2984 ( .IN(n1707), .OUT(n5221) );
  NAND2 U2985 ( .A(n5221), .B(n1706), .OUT(n4399) );
  NAND2 U2986 ( .A(n3247), .B(n4399), .OUT(n1817) );
  NAND2 U2987 ( .A(\mult_49/ab[11][18] ), .B(n1707), .OUT(n1816) );
  INV U2988 ( .IN(n1815), .OUT(n5222) );
  NAND2 U2989 ( .A(n5222), .B(n1814), .OUT(n4461) );
  NAND2 U2990 ( .A(n3328), .B(n4461), .OUT(n4835) );
  NAND2 U2991 ( .A(\mult_49/ab[12][18] ), .B(n1815), .OUT(n4462) );
  NAND2 U2992 ( .A(n5081), .B(n853), .OUT(n5223) );
  NAND2 U2993 ( .A(n2605), .B(n5223), .OUT(n921) );
  NAND2 U2994 ( .A(\mult_49/ab[2][17] ), .B(n850), .OUT(n920) );
  INV U2995 ( .IN(n919), .OUT(n5224) );
  NAND2 U2996 ( .A(n5224), .B(n918), .OUT(n4014) );
  NAND2 U2997 ( .A(n2656), .B(n4014), .OUT(n993) );
  NAND2 U2998 ( .A(\mult_49/ab[3][17] ), .B(n919), .OUT(n992) );
  INV U2999 ( .IN(n991), .OUT(n5225) );
  NAND2 U3000 ( .A(n5225), .B(n990), .OUT(n4049) );
  NAND2 U3001 ( .A(n2710), .B(n4049), .OUT(n1069) );
  NAND2 U3002 ( .A(\mult_49/ab[4][17] ), .B(n991), .OUT(n1068) );
  INV U3003 ( .IN(n1067), .OUT(n5226) );
  NAND2 U3004 ( .A(n5226), .B(n1066), .OUT(n4086) );
  NAND2 U3005 ( .A(n2767), .B(n4086), .OUT(n1149) );
  NAND2 U3006 ( .A(\mult_49/ab[5][17] ), .B(n1067), .OUT(n1148) );
  INV U3007 ( .IN(n1147), .OUT(n5227) );
  NAND2 U3008 ( .A(n5227), .B(n1146), .OUT(n4125) );
  NAND2 U3009 ( .A(n2827), .B(n4125), .OUT(n1233) );
  NAND2 U3010 ( .A(\mult_49/ab[6][17] ), .B(n1147), .OUT(n1232) );
  INV U3011 ( .IN(n1231), .OUT(n5228) );
  NAND2 U3012 ( .A(n5228), .B(n1230), .OUT(n4166) );
  NAND2 U3013 ( .A(n2890), .B(n4166), .OUT(n1321) );
  NAND2 U3014 ( .A(\mult_49/ab[7][17] ), .B(n1231), .OUT(n1320) );
  INV U3015 ( .IN(n1319), .OUT(n5229) );
  NAND2 U3016 ( .A(n5229), .B(n1318), .OUT(n4209) );
  NAND2 U3017 ( .A(n2956), .B(n4209), .OUT(n1413) );
  NAND2 U3018 ( .A(\mult_49/ab[8][17] ), .B(n1319), .OUT(n1412) );
  INV U3019 ( .IN(n1411), .OUT(n5230) );
  NAND2 U3020 ( .A(n5230), .B(n1410), .OUT(n4254) );
  NAND2 U3021 ( .A(n3025), .B(n4254), .OUT(n1509) );
  NAND2 U3022 ( .A(\mult_49/ab[9][17] ), .B(n1411), .OUT(n1508) );
  INV U3023 ( .IN(n1507), .OUT(n5231) );
  NAND2 U3024 ( .A(n5231), .B(n1506), .OUT(n4301) );
  NAND2 U3025 ( .A(n3097), .B(n4301), .OUT(n1609) );
  NAND2 U3026 ( .A(\mult_49/ab[10][17] ), .B(n1507), .OUT(n1608) );
  INV U3027 ( .IN(n1607), .OUT(n5232) );
  NAND2 U3028 ( .A(n5232), .B(n1606), .OUT(n4350) );
  NAND2 U3029 ( .A(n3172), .B(n4350), .OUT(n1713) );
  NAND2 U3030 ( .A(\mult_49/ab[11][17] ), .B(n1607), .OUT(n1712) );
  INV U3031 ( .IN(n1711), .OUT(n5233) );
  NAND2 U3032 ( .A(n5233), .B(n1710), .OUT(n4401) );
  NAND2 U3033 ( .A(n3250), .B(n4401), .OUT(n1821) );
  NAND2 U3034 ( .A(\mult_49/ab[12][17] ), .B(n1711), .OUT(n1820) );
  INV U3035 ( .IN(n1819), .OUT(n5234) );
  NAND2 U3036 ( .A(n5234), .B(n1818), .OUT(n4464) );
  NAND2 U3037 ( .A(n3331), .B(n4464), .OUT(n4805) );
  NAND2 U3038 ( .A(\mult_49/ab[13][17] ), .B(n1819), .OUT(n4465) );
  NAND2 U3039 ( .A(n5082), .B(n793), .OUT(n5235) );
  NAND2 U3040 ( .A(n2560), .B(n5235), .OUT(n857) );
  NAND2 U3041 ( .A(\mult_49/ab[2][16] ), .B(n790), .OUT(n856) );
  INV U3042 ( .IN(n855), .OUT(n5236) );
  NAND2 U3043 ( .A(n5236), .B(n854), .OUT(n3983) );
  NAND2 U3044 ( .A(n2608), .B(n3983), .OUT(n925) );
  NAND2 U3045 ( .A(\mult_49/ab[3][16] ), .B(n855), .OUT(n924) );
  INV U3046 ( .IN(n923), .OUT(n5237) );
  NAND2 U3047 ( .A(n5237), .B(n922), .OUT(n4016) );
  NAND2 U3048 ( .A(n2659), .B(n4016), .OUT(n997) );
  NAND2 U3049 ( .A(\mult_49/ab[4][16] ), .B(n923), .OUT(n996) );
  INV U3050 ( .IN(n995), .OUT(n5238) );
  NAND2 U3051 ( .A(n5238), .B(n994), .OUT(n4051) );
  NAND2 U3052 ( .A(n2713), .B(n4051), .OUT(n1073) );
  NAND2 U3053 ( .A(\mult_49/ab[5][16] ), .B(n995), .OUT(n1072) );
  INV U3054 ( .IN(n1071), .OUT(n5239) );
  NAND2 U3055 ( .A(n5239), .B(n1070), .OUT(n4088) );
  NAND2 U3056 ( .A(n2770), .B(n4088), .OUT(n1153) );
  NAND2 U3057 ( .A(\mult_49/ab[6][16] ), .B(n1071), .OUT(n1152) );
  INV U3058 ( .IN(n1151), .OUT(n5240) );
  NAND2 U3059 ( .A(n5240), .B(n1150), .OUT(n4127) );
  NAND2 U3060 ( .A(n2830), .B(n4127), .OUT(n1237) );
  NAND2 U3061 ( .A(\mult_49/ab[7][16] ), .B(n1151), .OUT(n1236) );
  INV U3062 ( .IN(n1235), .OUT(n5241) );
  NAND2 U3063 ( .A(n5241), .B(n1234), .OUT(n4168) );
  NAND2 U3064 ( .A(n2893), .B(n4168), .OUT(n1325) );
  NAND2 U3065 ( .A(\mult_49/ab[8][16] ), .B(n1235), .OUT(n1324) );
  INV U3066 ( .IN(n1323), .OUT(n5242) );
  NAND2 U3067 ( .A(n5242), .B(n1322), .OUT(n4211) );
  NAND2 U3068 ( .A(n2959), .B(n4211), .OUT(n1417) );
  NAND2 U3069 ( .A(\mult_49/ab[9][16] ), .B(n1323), .OUT(n1416) );
  INV U3070 ( .IN(n1415), .OUT(n5243) );
  NAND2 U3071 ( .A(n5243), .B(n1414), .OUT(n4256) );
  NAND2 U3072 ( .A(n3028), .B(n4256), .OUT(n1513) );
  NAND2 U3073 ( .A(\mult_49/ab[10][16] ), .B(n1415), .OUT(n1512) );
  INV U3074 ( .IN(n1511), .OUT(n5244) );
  NAND2 U3075 ( .A(n5244), .B(n1510), .OUT(n4303) );
  NAND2 U3076 ( .A(n3100), .B(n4303), .OUT(n1613) );
  NAND2 U3077 ( .A(\mult_49/ab[11][16] ), .B(n1511), .OUT(n1612) );
  INV U3078 ( .IN(n1611), .OUT(n5245) );
  NAND2 U3079 ( .A(n5245), .B(n1610), .OUT(n4352) );
  NAND2 U3080 ( .A(n3175), .B(n4352), .OUT(n1717) );
  NAND2 U3081 ( .A(\mult_49/ab[12][16] ), .B(n1611), .OUT(n1716) );
  INV U3082 ( .IN(n1715), .OUT(n5246) );
  NAND2 U3083 ( .A(n5246), .B(n1714), .OUT(n4403) );
  NAND2 U3084 ( .A(n3253), .B(n4403), .OUT(n1825) );
  NAND2 U3085 ( .A(\mult_49/ab[13][16] ), .B(n1715), .OUT(n1824) );
  INV U3086 ( .IN(n1823), .OUT(n5247) );
  NAND2 U3087 ( .A(n5247), .B(n1822), .OUT(n4467) );
  NAND2 U3088 ( .A(n3334), .B(n4467), .OUT(n4807) );
  NAND2 U3089 ( .A(\mult_49/ab[14][16] ), .B(n1823), .OUT(n4468) );
  NAND2 U3090 ( .A(n5083), .B(n737), .OUT(n5248) );
  NAND2 U3091 ( .A(n2518), .B(n5248), .OUT(n797) );
  NAND2 U3092 ( .A(\mult_49/ab[2][15] ), .B(n734), .OUT(n796) );
  INV U3093 ( .IN(n795), .OUT(n5249) );
  NAND2 U3094 ( .A(n5249), .B(n794), .OUT(n3954) );
  NAND2 U3095 ( .A(n2563), .B(n3954), .OUT(n861) );
  NAND2 U3096 ( .A(\mult_49/ab[3][15] ), .B(n795), .OUT(n860) );
  INV U3097 ( .IN(n859), .OUT(n5250) );
  NAND2 U3098 ( .A(n5250), .B(n858), .OUT(n3985) );
  NAND2 U3099 ( .A(n2611), .B(n3985), .OUT(n929) );
  NAND2 U3100 ( .A(\mult_49/ab[4][15] ), .B(n859), .OUT(n928) );
  INV U3101 ( .IN(n927), .OUT(n5251) );
  NAND2 U3102 ( .A(n5251), .B(n926), .OUT(n4018) );
  NAND2 U3103 ( .A(n2662), .B(n4018), .OUT(n1001) );
  NAND2 U3104 ( .A(\mult_49/ab[5][15] ), .B(n927), .OUT(n1000) );
  INV U3105 ( .IN(n999), .OUT(n5252) );
  NAND2 U3106 ( .A(n5252), .B(n998), .OUT(n4053) );
  NAND2 U3107 ( .A(n2716), .B(n4053), .OUT(n1077) );
  NAND2 U3108 ( .A(\mult_49/ab[6][15] ), .B(n999), .OUT(n1076) );
  INV U3109 ( .IN(n1075), .OUT(n5253) );
  NAND2 U3110 ( .A(n5253), .B(n1074), .OUT(n4090) );
  NAND2 U3111 ( .A(n2773), .B(n4090), .OUT(n1157) );
  NAND2 U3112 ( .A(\mult_49/ab[7][15] ), .B(n1075), .OUT(n1156) );
  INV U3113 ( .IN(n1155), .OUT(n5254) );
  NAND2 U3114 ( .A(n5254), .B(n1154), .OUT(n4129) );
  NAND2 U3115 ( .A(n2833), .B(n4129), .OUT(n1241) );
  NAND2 U3116 ( .A(\mult_49/ab[8][15] ), .B(n1155), .OUT(n1240) );
  INV U3117 ( .IN(n1239), .OUT(n5255) );
  NAND2 U3118 ( .A(n5255), .B(n1238), .OUT(n4170) );
  NAND2 U3119 ( .A(n2896), .B(n4170), .OUT(n1329) );
  NAND2 U3120 ( .A(\mult_49/ab[9][15] ), .B(n1239), .OUT(n1328) );
  INV U3121 ( .IN(n1327), .OUT(n5256) );
  NAND2 U3122 ( .A(n5256), .B(n1326), .OUT(n4213) );
  NAND2 U3123 ( .A(n2962), .B(n4213), .OUT(n1421) );
  NAND2 U3124 ( .A(\mult_49/ab[10][15] ), .B(n1327), .OUT(n1420) );
  INV U3125 ( .IN(n1419), .OUT(n5257) );
  NAND2 U3126 ( .A(n5257), .B(n1418), .OUT(n4258) );
  NAND2 U3127 ( .A(n3031), .B(n4258), .OUT(n1517) );
  NAND2 U3128 ( .A(\mult_49/ab[11][15] ), .B(n1419), .OUT(n1516) );
  INV U3129 ( .IN(n1515), .OUT(n5258) );
  NAND2 U3130 ( .A(n5258), .B(n1514), .OUT(n4305) );
  NAND2 U3131 ( .A(n3103), .B(n4305), .OUT(n1617) );
  NAND2 U3132 ( .A(\mult_49/ab[12][15] ), .B(n1515), .OUT(n1616) );
  INV U3133 ( .IN(n1615), .OUT(n5259) );
  NAND2 U3134 ( .A(n5259), .B(n1614), .OUT(n4354) );
  NAND2 U3135 ( .A(n3178), .B(n4354), .OUT(n1721) );
  NAND2 U3136 ( .A(\mult_49/ab[13][15] ), .B(n1615), .OUT(n1720) );
  INV U3137 ( .IN(n1719), .OUT(n5260) );
  NAND2 U3138 ( .A(n5260), .B(n1718), .OUT(n4405) );
  NAND2 U3139 ( .A(n3256), .B(n4405), .OUT(n1829) );
  NAND2 U3140 ( .A(\mult_49/ab[14][15] ), .B(n1719), .OUT(n1828) );
  INV U3141 ( .IN(n1827), .OUT(n5261) );
  NAND2 U3142 ( .A(n5261), .B(n1826), .OUT(n4470) );
  NAND2 U3143 ( .A(n3337), .B(n4470), .OUT(n4811) );
  NAND2 U3144 ( .A(\mult_49/ab[15][15] ), .B(n1827), .OUT(n4471) );
  NAND2 U3145 ( .A(n5084), .B(n685), .OUT(n5262) );
  NAND2 U3146 ( .A(n2479), .B(n5262), .OUT(n741) );
  NAND2 U3147 ( .A(\mult_49/ab[2][14] ), .B(n682), .OUT(n740) );
  INV U3148 ( .IN(n739), .OUT(n5263) );
  NAND2 U3149 ( .A(n5263), .B(n738), .OUT(n3927) );
  NAND2 U3150 ( .A(n2521), .B(n3927), .OUT(n801) );
  NAND2 U3151 ( .A(\mult_49/ab[3][14] ), .B(n739), .OUT(n800) );
  INV U3152 ( .IN(n799), .OUT(n5264) );
  NAND2 U3153 ( .A(n5264), .B(n798), .OUT(n3956) );
  NAND2 U3154 ( .A(n2566), .B(n3956), .OUT(n865) );
  NAND2 U3155 ( .A(\mult_49/ab[4][14] ), .B(n799), .OUT(n864) );
  INV U3156 ( .IN(n863), .OUT(n5265) );
  NAND2 U3157 ( .A(n5265), .B(n862), .OUT(n3987) );
  NAND2 U3158 ( .A(n2614), .B(n3987), .OUT(n933) );
  NAND2 U3159 ( .A(\mult_49/ab[5][14] ), .B(n863), .OUT(n932) );
  INV U3160 ( .IN(n931), .OUT(n5266) );
  NAND2 U3161 ( .A(n5266), .B(n930), .OUT(n4020) );
  NAND2 U3162 ( .A(n2665), .B(n4020), .OUT(n1005) );
  NAND2 U3163 ( .A(\mult_49/ab[6][14] ), .B(n931), .OUT(n1004) );
  INV U3164 ( .IN(n1003), .OUT(n5267) );
  NAND2 U3165 ( .A(n5267), .B(n1002), .OUT(n4055) );
  NAND2 U3166 ( .A(n2719), .B(n4055), .OUT(n1081) );
  NAND2 U3167 ( .A(\mult_49/ab[7][14] ), .B(n1003), .OUT(n1080) );
  INV U3168 ( .IN(n1079), .OUT(n5268) );
  NAND2 U3169 ( .A(n5268), .B(n1078), .OUT(n4092) );
  NAND2 U3170 ( .A(n2776), .B(n4092), .OUT(n1161) );
  NAND2 U3171 ( .A(\mult_49/ab[8][14] ), .B(n1079), .OUT(n1160) );
  INV U3172 ( .IN(n1159), .OUT(n5269) );
  NAND2 U3173 ( .A(n5269), .B(n1158), .OUT(n4131) );
  NAND2 U3174 ( .A(n2836), .B(n4131), .OUT(n1245) );
  NAND2 U3175 ( .A(\mult_49/ab[9][14] ), .B(n1159), .OUT(n1244) );
  INV U3176 ( .IN(n1243), .OUT(n5270) );
  NAND2 U3177 ( .A(n5270), .B(n1242), .OUT(n4172) );
  NAND2 U3178 ( .A(n2899), .B(n4172), .OUT(n1333) );
  NAND2 U3179 ( .A(\mult_49/ab[10][14] ), .B(n1243), .OUT(n1332) );
  INV U3180 ( .IN(n1331), .OUT(n5271) );
  NAND2 U3181 ( .A(n5271), .B(n1330), .OUT(n4215) );
  NAND2 U3182 ( .A(n2965), .B(n4215), .OUT(n1425) );
  NAND2 U3183 ( .A(\mult_49/ab[11][14] ), .B(n1331), .OUT(n1424) );
  INV U3184 ( .IN(n1423), .OUT(n5272) );
  NAND2 U3185 ( .A(n5272), .B(n1422), .OUT(n4260) );
  NAND2 U3186 ( .A(n3034), .B(n4260), .OUT(n1521) );
  NAND2 U3187 ( .A(\mult_49/ab[12][14] ), .B(n1423), .OUT(n1520) );
  INV U3188 ( .IN(n1519), .OUT(n5273) );
  NAND2 U3189 ( .A(n5273), .B(n1518), .OUT(n4307) );
  NAND2 U3190 ( .A(n3106), .B(n4307), .OUT(n1621) );
  NAND2 U3191 ( .A(\mult_49/ab[13][14] ), .B(n1519), .OUT(n1620) );
  INV U3192 ( .IN(n1619), .OUT(n5274) );
  NAND2 U3193 ( .A(n5274), .B(n1618), .OUT(n4356) );
  NAND2 U3194 ( .A(n3181), .B(n4356), .OUT(n1725) );
  NAND2 U3195 ( .A(\mult_49/ab[14][14] ), .B(n1619), .OUT(n1724) );
  INV U3196 ( .IN(n1723), .OUT(n5275) );
  NAND2 U3197 ( .A(n5275), .B(n1722), .OUT(n4407) );
  NAND2 U3198 ( .A(n3259), .B(n4407), .OUT(n1833) );
  NAND2 U3199 ( .A(\mult_49/ab[15][14] ), .B(n1723), .OUT(n1832) );
  INV U3200 ( .IN(n1831), .OUT(n5276) );
  NAND2 U3201 ( .A(n5276), .B(n1830), .OUT(n4473) );
  NAND2 U3202 ( .A(n3340), .B(n4473), .OUT(n4799) );
  NAND2 U3203 ( .A(\mult_49/ab[16][14] ), .B(n1831), .OUT(n4474) );
  NAND2 U3204 ( .A(n5085), .B(n637), .OUT(n5277) );
  NAND2 U3205 ( .A(n2443), .B(n5277), .OUT(n689) );
  NAND2 U3206 ( .A(\mult_49/ab[2][13] ), .B(n634), .OUT(n688) );
  INV U3207 ( .IN(n687), .OUT(n5278) );
  NAND2 U3208 ( .A(n5278), .B(n686), .OUT(n3902) );
  NAND2 U3209 ( .A(n2482), .B(n3902), .OUT(n745) );
  NAND2 U3210 ( .A(\mult_49/ab[3][13] ), .B(n687), .OUT(n744) );
  INV U3211 ( .IN(n743), .OUT(n5279) );
  NAND2 U3212 ( .A(n5279), .B(n742), .OUT(n3929) );
  NAND2 U3213 ( .A(n2524), .B(n3929), .OUT(n805) );
  NAND2 U3214 ( .A(\mult_49/ab[4][13] ), .B(n743), .OUT(n804) );
  INV U3215 ( .IN(n803), .OUT(n5280) );
  NAND2 U3216 ( .A(n5280), .B(n802), .OUT(n3958) );
  NAND2 U3217 ( .A(n2569), .B(n3958), .OUT(n869) );
  NAND2 U3218 ( .A(\mult_49/ab[5][13] ), .B(n803), .OUT(n868) );
  INV U3219 ( .IN(n867), .OUT(n5281) );
  NAND2 U3220 ( .A(n5281), .B(n866), .OUT(n3989) );
  NAND2 U3221 ( .A(n2617), .B(n3989), .OUT(n937) );
  NAND2 U3222 ( .A(\mult_49/ab[6][13] ), .B(n867), .OUT(n936) );
  INV U3223 ( .IN(n935), .OUT(n5282) );
  NAND2 U3224 ( .A(n5282), .B(n934), .OUT(n4022) );
  NAND2 U3225 ( .A(n2668), .B(n4022), .OUT(n1009) );
  NAND2 U3226 ( .A(\mult_49/ab[7][13] ), .B(n935), .OUT(n1008) );
  INV U3227 ( .IN(n1007), .OUT(n5283) );
  NAND2 U3228 ( .A(n5283), .B(n1006), .OUT(n4057) );
  NAND2 U3229 ( .A(n2722), .B(n4057), .OUT(n1085) );
  NAND2 U3230 ( .A(\mult_49/ab[8][13] ), .B(n1007), .OUT(n1084) );
  INV U3231 ( .IN(n1083), .OUT(n5284) );
  NAND2 U3232 ( .A(n5284), .B(n1082), .OUT(n4094) );
  NAND2 U3233 ( .A(n2779), .B(n4094), .OUT(n1165) );
  NAND2 U3234 ( .A(\mult_49/ab[9][13] ), .B(n1083), .OUT(n1164) );
  INV U3235 ( .IN(n1163), .OUT(n5285) );
  NAND2 U3236 ( .A(n5285), .B(n1162), .OUT(n4133) );
  NAND2 U3237 ( .A(n2839), .B(n4133), .OUT(n1249) );
  NAND2 U3238 ( .A(\mult_49/ab[10][13] ), .B(n1163), .OUT(n1248) );
  INV U3239 ( .IN(n1247), .OUT(n5286) );
  NAND2 U3240 ( .A(n5286), .B(n1246), .OUT(n4174) );
  NAND2 U3241 ( .A(n2902), .B(n4174), .OUT(n1337) );
  NAND2 U3242 ( .A(\mult_49/ab[11][13] ), .B(n1247), .OUT(n1336) );
  INV U3243 ( .IN(n1335), .OUT(n5287) );
  NAND2 U3244 ( .A(n5287), .B(n1334), .OUT(n4217) );
  NAND2 U3245 ( .A(n2968), .B(n4217), .OUT(n1429) );
  NAND2 U3246 ( .A(\mult_49/ab[12][13] ), .B(n1335), .OUT(n1428) );
  INV U3247 ( .IN(n1427), .OUT(n5288) );
  NAND2 U3248 ( .A(n5288), .B(n1426), .OUT(n4262) );
  NAND2 U3249 ( .A(n3037), .B(n4262), .OUT(n1525) );
  NAND2 U3250 ( .A(\mult_49/ab[13][13] ), .B(n1427), .OUT(n1524) );
  INV U3251 ( .IN(n1523), .OUT(n5289) );
  NAND2 U3252 ( .A(n5289), .B(n1522), .OUT(n4309) );
  NAND2 U3253 ( .A(n3109), .B(n4309), .OUT(n1625) );
  NAND2 U3254 ( .A(\mult_49/ab[14][13] ), .B(n1523), .OUT(n1624) );
  INV U3255 ( .IN(n1623), .OUT(n5290) );
  NAND2 U3256 ( .A(n5290), .B(n1622), .OUT(n4358) );
  NAND2 U3257 ( .A(n3184), .B(n4358), .OUT(n1729) );
  NAND2 U3258 ( .A(\mult_49/ab[15][13] ), .B(n1623), .OUT(n1728) );
  INV U3259 ( .IN(n1727), .OUT(n5291) );
  NAND2 U3260 ( .A(n5291), .B(n1726), .OUT(n4409) );
  NAND2 U3261 ( .A(n3262), .B(n4409), .OUT(n1837) );
  NAND2 U3262 ( .A(\mult_49/ab[16][13] ), .B(n1727), .OUT(n1836) );
  INV U3263 ( .IN(n1835), .OUT(n5292) );
  NAND2 U3264 ( .A(n5292), .B(n1834), .OUT(n4476) );
  NAND2 U3265 ( .A(n3343), .B(n4476), .OUT(n4837) );
  NAND2 U3266 ( .A(\mult_49/ab[17][13] ), .B(n1835), .OUT(n4477) );
  NAND2 U3267 ( .A(n5086), .B(n593), .OUT(n5293) );
  NAND2 U3268 ( .A(n2410), .B(n5293), .OUT(n641) );
  NAND2 U3269 ( .A(\mult_49/ab[2][12] ), .B(n590), .OUT(n640) );
  INV U3270 ( .IN(n639), .OUT(n5294) );
  NAND2 U3271 ( .A(n5294), .B(n638), .OUT(n3879) );
  NAND2 U3272 ( .A(n2446), .B(n3879), .OUT(n693) );
  NAND2 U3273 ( .A(\mult_49/ab[3][12] ), .B(n639), .OUT(n692) );
  INV U3274 ( .IN(n691), .OUT(n5295) );
  NAND2 U3275 ( .A(n5295), .B(n690), .OUT(n3904) );
  NAND2 U3276 ( .A(n2485), .B(n3904), .OUT(n749) );
  NAND2 U3277 ( .A(\mult_49/ab[4][12] ), .B(n691), .OUT(n748) );
  INV U3278 ( .IN(n747), .OUT(n5296) );
  NAND2 U3279 ( .A(n5296), .B(n746), .OUT(n3931) );
  NAND2 U3280 ( .A(n2527), .B(n3931), .OUT(n809) );
  NAND2 U3281 ( .A(\mult_49/ab[5][12] ), .B(n747), .OUT(n808) );
  INV U3282 ( .IN(n807), .OUT(n5297) );
  NAND2 U3283 ( .A(n5297), .B(n806), .OUT(n3960) );
  NAND2 U3284 ( .A(n2572), .B(n3960), .OUT(n873) );
  NAND2 U3285 ( .A(\mult_49/ab[6][12] ), .B(n807), .OUT(n872) );
  INV U3286 ( .IN(n871), .OUT(n5298) );
  NAND2 U3287 ( .A(n5298), .B(n870), .OUT(n3991) );
  NAND2 U3288 ( .A(n2620), .B(n3991), .OUT(n941) );
  NAND2 U3289 ( .A(\mult_49/ab[7][12] ), .B(n871), .OUT(n940) );
  INV U3290 ( .IN(n939), .OUT(n5299) );
  NAND2 U3291 ( .A(n5299), .B(n938), .OUT(n4024) );
  NAND2 U3292 ( .A(n2671), .B(n4024), .OUT(n1013) );
  NAND2 U3293 ( .A(\mult_49/ab[8][12] ), .B(n939), .OUT(n1012) );
  INV U3294 ( .IN(n1011), .OUT(n5300) );
  NAND2 U3295 ( .A(n5300), .B(n1010), .OUT(n4059) );
  NAND2 U3296 ( .A(n2725), .B(n4059), .OUT(n1089) );
  NAND2 U3297 ( .A(\mult_49/ab[9][12] ), .B(n1011), .OUT(n1088) );
  INV U3298 ( .IN(n1087), .OUT(n5301) );
  NAND2 U3299 ( .A(n5301), .B(n1086), .OUT(n4096) );
  NAND2 U3300 ( .A(n2782), .B(n4096), .OUT(n1169) );
  NAND2 U3301 ( .A(\mult_49/ab[10][12] ), .B(n1087), .OUT(n1168) );
  INV U3302 ( .IN(n1167), .OUT(n5302) );
  NAND2 U3303 ( .A(n5302), .B(n1166), .OUT(n4135) );
  NAND2 U3304 ( .A(n2842), .B(n4135), .OUT(n1253) );
  NAND2 U3305 ( .A(\mult_49/ab[11][12] ), .B(n1167), .OUT(n1252) );
  INV U3306 ( .IN(n1251), .OUT(n5303) );
  NAND2 U3307 ( .A(n5303), .B(n1250), .OUT(n4176) );
  NAND2 U3308 ( .A(n2905), .B(n4176), .OUT(n1341) );
  NAND2 U3309 ( .A(\mult_49/ab[12][12] ), .B(n1251), .OUT(n1340) );
  INV U3310 ( .IN(n1339), .OUT(n5304) );
  NAND2 U3311 ( .A(n5304), .B(n1338), .OUT(n4219) );
  NAND2 U3312 ( .A(n2971), .B(n4219), .OUT(n1433) );
  NAND2 U3313 ( .A(\mult_49/ab[13][12] ), .B(n1339), .OUT(n1432) );
  INV U3314 ( .IN(n1431), .OUT(n5305) );
  NAND2 U3315 ( .A(n5305), .B(n1430), .OUT(n4264) );
  NAND2 U3316 ( .A(n3040), .B(n4264), .OUT(n1529) );
  NAND2 U3317 ( .A(\mult_49/ab[14][12] ), .B(n1431), .OUT(n1528) );
  INV U3318 ( .IN(n1527), .OUT(n5306) );
  NAND2 U3319 ( .A(n5306), .B(n1526), .OUT(n4311) );
  NAND2 U3320 ( .A(n3112), .B(n4311), .OUT(n1629) );
  NAND2 U3321 ( .A(\mult_49/ab[15][12] ), .B(n1527), .OUT(n1628) );
  INV U3322 ( .IN(n1627), .OUT(n5307) );
  NAND2 U3323 ( .A(n5307), .B(n1626), .OUT(n4360) );
  NAND2 U3324 ( .A(n3187), .B(n4360), .OUT(n1733) );
  NAND2 U3325 ( .A(\mult_49/ab[16][12] ), .B(n1627), .OUT(n1732) );
  INV U3326 ( .IN(n1731), .OUT(n5308) );
  NAND2 U3327 ( .A(n5308), .B(n1730), .OUT(n4411) );
  NAND2 U3328 ( .A(n3265), .B(n4411), .OUT(n1841) );
  NAND2 U3329 ( .A(\mult_49/ab[17][12] ), .B(n1731), .OUT(n1840) );
  INV U3330 ( .IN(n1839), .OUT(n5309) );
  NAND2 U3331 ( .A(n5309), .B(n1838), .OUT(n4479) );
  NAND2 U3332 ( .A(n3346), .B(n4479), .OUT(n4839) );
  NAND2 U3333 ( .A(\mult_49/ab[18][12] ), .B(n1839), .OUT(n4480) );
  NAND2 U3334 ( .A(n5087), .B(n553), .OUT(n5310) );
  NAND2 U3335 ( .A(n2380), .B(n5310), .OUT(n597) );
  NAND2 U3336 ( .A(\mult_49/ab[2][11] ), .B(n550), .OUT(n596) );
  INV U3337 ( .IN(n595), .OUT(n5311) );
  NAND2 U3338 ( .A(n5311), .B(n594), .OUT(n3858) );
  NAND2 U3339 ( .A(n2413), .B(n3858), .OUT(n645) );
  NAND2 U3340 ( .A(\mult_49/ab[3][11] ), .B(n595), .OUT(n644) );
  INV U3341 ( .IN(n643), .OUT(n5312) );
  NAND2 U3342 ( .A(n5312), .B(n642), .OUT(n3881) );
  NAND2 U3343 ( .A(n2449), .B(n3881), .OUT(n697) );
  NAND2 U3344 ( .A(\mult_49/ab[4][11] ), .B(n643), .OUT(n696) );
  INV U3345 ( .IN(n695), .OUT(n5313) );
  NAND2 U3346 ( .A(n5313), .B(n694), .OUT(n3906) );
  NAND2 U3347 ( .A(n2488), .B(n3906), .OUT(n753) );
  NAND2 U3348 ( .A(\mult_49/ab[5][11] ), .B(n695), .OUT(n752) );
  INV U3349 ( .IN(n751), .OUT(n5314) );
  NAND2 U3350 ( .A(n5314), .B(n750), .OUT(n3933) );
  NAND2 U3351 ( .A(n2530), .B(n3933), .OUT(n813) );
  NAND2 U3352 ( .A(\mult_49/ab[6][11] ), .B(n751), .OUT(n812) );
  INV U3353 ( .IN(n811), .OUT(n5315) );
  NAND2 U3354 ( .A(n5315), .B(n810), .OUT(n3962) );
  NAND2 U3355 ( .A(n2575), .B(n3962), .OUT(n877) );
  NAND2 U3356 ( .A(\mult_49/ab[7][11] ), .B(n811), .OUT(n876) );
  INV U3357 ( .IN(n875), .OUT(n5316) );
  NAND2 U3358 ( .A(n5316), .B(n874), .OUT(n3993) );
  NAND2 U3359 ( .A(n2623), .B(n3993), .OUT(n945) );
  NAND2 U3360 ( .A(\mult_49/ab[8][11] ), .B(n875), .OUT(n944) );
  INV U3361 ( .IN(n943), .OUT(n5317) );
  NAND2 U3362 ( .A(n5317), .B(n942), .OUT(n4026) );
  NAND2 U3363 ( .A(n2674), .B(n4026), .OUT(n1017) );
  NAND2 U3364 ( .A(\mult_49/ab[9][11] ), .B(n943), .OUT(n1016) );
  INV U3365 ( .IN(n1015), .OUT(n5318) );
  NAND2 U3366 ( .A(n5318), .B(n1014), .OUT(n4061) );
  NAND2 U3367 ( .A(n2728), .B(n4061), .OUT(n1093) );
  NAND2 U3368 ( .A(\mult_49/ab[10][11] ), .B(n1015), .OUT(n1092) );
  INV U3369 ( .IN(n1091), .OUT(n5319) );
  NAND2 U3370 ( .A(n5319), .B(n1090), .OUT(n4098) );
  NAND2 U3371 ( .A(n2785), .B(n4098), .OUT(n1173) );
  NAND2 U3372 ( .A(\mult_49/ab[11][11] ), .B(n1091), .OUT(n1172) );
  INV U3373 ( .IN(n1171), .OUT(n5320) );
  NAND2 U3374 ( .A(n5320), .B(n1170), .OUT(n4137) );
  NAND2 U3375 ( .A(n2845), .B(n4137), .OUT(n1257) );
  NAND2 U3376 ( .A(\mult_49/ab[12][11] ), .B(n1171), .OUT(n1256) );
  INV U3377 ( .IN(n1255), .OUT(n5321) );
  NAND2 U3378 ( .A(n5321), .B(n1254), .OUT(n4178) );
  NAND2 U3379 ( .A(n2908), .B(n4178), .OUT(n1345) );
  NAND2 U3380 ( .A(\mult_49/ab[13][11] ), .B(n1255), .OUT(n1344) );
  INV U3381 ( .IN(n1343), .OUT(n5322) );
  NAND2 U3382 ( .A(n5322), .B(n1342), .OUT(n4221) );
  NAND2 U3383 ( .A(n2974), .B(n4221), .OUT(n1437) );
  NAND2 U3384 ( .A(\mult_49/ab[14][11] ), .B(n1343), .OUT(n1436) );
  INV U3385 ( .IN(n1435), .OUT(n5323) );
  NAND2 U3386 ( .A(n5323), .B(n1434), .OUT(n4266) );
  NAND2 U3387 ( .A(n3043), .B(n4266), .OUT(n1533) );
  NAND2 U3388 ( .A(\mult_49/ab[15][11] ), .B(n1435), .OUT(n1532) );
  INV U3389 ( .IN(n1531), .OUT(n5324) );
  NAND2 U3390 ( .A(n5324), .B(n1530), .OUT(n4313) );
  NAND2 U3391 ( .A(n3115), .B(n4313), .OUT(n1633) );
  NAND2 U3392 ( .A(\mult_49/ab[16][11] ), .B(n1531), .OUT(n1632) );
  INV U3393 ( .IN(n1631), .OUT(n5325) );
  NAND2 U3394 ( .A(n5325), .B(n1630), .OUT(n4362) );
  NAND2 U3395 ( .A(n3190), .B(n4362), .OUT(n1737) );
  NAND2 U3396 ( .A(\mult_49/ab[17][11] ), .B(n1631), .OUT(n1736) );
  INV U3397 ( .IN(n1735), .OUT(n5326) );
  NAND2 U3398 ( .A(n5326), .B(n1734), .OUT(n4413) );
  NAND2 U3399 ( .A(n3268), .B(n4413), .OUT(n1845) );
  NAND2 U3400 ( .A(\mult_49/ab[18][11] ), .B(n1735), .OUT(n1844) );
  INV U3401 ( .IN(n1843), .OUT(n5327) );
  NAND2 U3402 ( .A(n5327), .B(n1842), .OUT(n4482) );
  NAND2 U3403 ( .A(n3349), .B(n4482), .OUT(n4813) );
  NAND2 U3404 ( .A(\mult_49/ab[19][11] ), .B(n1843), .OUT(n4483) );
  NAND2 U3405 ( .A(n5088), .B(n517), .OUT(n5328) );
  NAND2 U3406 ( .A(n2353), .B(n5328), .OUT(n557) );
  NAND2 U3407 ( .A(\mult_49/ab[2][10] ), .B(n514), .OUT(n556) );
  INV U3408 ( .IN(n555), .OUT(n5329) );
  NAND2 U3409 ( .A(n5329), .B(n554), .OUT(n3839) );
  NAND2 U3410 ( .A(n2383), .B(n3839), .OUT(n601) );
  NAND2 U3411 ( .A(\mult_49/ab[3][10] ), .B(n555), .OUT(n600) );
  INV U3412 ( .IN(n599), .OUT(n5330) );
  NAND2 U3413 ( .A(n5330), .B(n598), .OUT(n3860) );
  NAND2 U3414 ( .A(n2416), .B(n3860), .OUT(n649) );
  NAND2 U3415 ( .A(\mult_49/ab[4][10] ), .B(n599), .OUT(n648) );
  INV U3416 ( .IN(n647), .OUT(n5331) );
  NAND2 U3417 ( .A(n5331), .B(n646), .OUT(n3883) );
  NAND2 U3418 ( .A(n2452), .B(n3883), .OUT(n701) );
  NAND2 U3419 ( .A(\mult_49/ab[5][10] ), .B(n647), .OUT(n700) );
  INV U3420 ( .IN(n699), .OUT(n5332) );
  NAND2 U3421 ( .A(n5332), .B(n698), .OUT(n3908) );
  NAND2 U3422 ( .A(n2491), .B(n3908), .OUT(n757) );
  NAND2 U3423 ( .A(\mult_49/ab[6][10] ), .B(n699), .OUT(n756) );
  INV U3424 ( .IN(n755), .OUT(n5333) );
  NAND2 U3425 ( .A(n5333), .B(n754), .OUT(n3935) );
  NAND2 U3426 ( .A(n2533), .B(n3935), .OUT(n817) );
  NAND2 U3427 ( .A(\mult_49/ab[7][10] ), .B(n755), .OUT(n816) );
  INV U3428 ( .IN(n815), .OUT(n5334) );
  NAND2 U3429 ( .A(n5334), .B(n814), .OUT(n3964) );
  NAND2 U3430 ( .A(n2578), .B(n3964), .OUT(n881) );
  NAND2 U3431 ( .A(\mult_49/ab[8][10] ), .B(n815), .OUT(n880) );
  INV U3432 ( .IN(n879), .OUT(n5335) );
  NAND2 U3433 ( .A(n5335), .B(n878), .OUT(n3995) );
  NAND2 U3434 ( .A(n2626), .B(n3995), .OUT(n949) );
  NAND2 U3435 ( .A(\mult_49/ab[9][10] ), .B(n879), .OUT(n948) );
  INV U3436 ( .IN(n947), .OUT(n5336) );
  NAND2 U3437 ( .A(n5336), .B(n946), .OUT(n4028) );
  NAND2 U3438 ( .A(n2677), .B(n4028), .OUT(n1021) );
  NAND2 U3439 ( .A(\mult_49/ab[10][10] ), .B(n947), .OUT(n1020) );
  INV U3440 ( .IN(n1019), .OUT(n5337) );
  NAND2 U3441 ( .A(n5337), .B(n1018), .OUT(n4063) );
  NAND2 U3442 ( .A(n2731), .B(n4063), .OUT(n1097) );
  NAND2 U3443 ( .A(\mult_49/ab[11][10] ), .B(n1019), .OUT(n1096) );
  INV U3444 ( .IN(n1095), .OUT(n5338) );
  NAND2 U3445 ( .A(n5338), .B(n1094), .OUT(n4100) );
  NAND2 U3446 ( .A(n2788), .B(n4100), .OUT(n1177) );
  NAND2 U3447 ( .A(\mult_49/ab[12][10] ), .B(n1095), .OUT(n1176) );
  INV U3448 ( .IN(n1175), .OUT(n5339) );
  NAND2 U3449 ( .A(n5339), .B(n1174), .OUT(n4139) );
  NAND2 U3450 ( .A(n2848), .B(n4139), .OUT(n1261) );
  NAND2 U3451 ( .A(\mult_49/ab[13][10] ), .B(n1175), .OUT(n1260) );
  INV U3452 ( .IN(n1259), .OUT(n5340) );
  NAND2 U3453 ( .A(n5340), .B(n1258), .OUT(n4180) );
  NAND2 U3454 ( .A(n2911), .B(n4180), .OUT(n1349) );
  NAND2 U3455 ( .A(\mult_49/ab[14][10] ), .B(n1259), .OUT(n1348) );
  INV U3456 ( .IN(n1347), .OUT(n5341) );
  NAND2 U3457 ( .A(n5341), .B(n1346), .OUT(n4223) );
  NAND2 U3458 ( .A(n2977), .B(n4223), .OUT(n1441) );
  NAND2 U3459 ( .A(\mult_49/ab[15][10] ), .B(n1347), .OUT(n1440) );
  INV U3460 ( .IN(n1439), .OUT(n5342) );
  NAND2 U3461 ( .A(n5342), .B(n1438), .OUT(n4268) );
  NAND2 U3462 ( .A(n3046), .B(n4268), .OUT(n1537) );
  NAND2 U3463 ( .A(\mult_49/ab[16][10] ), .B(n1439), .OUT(n1536) );
  INV U3464 ( .IN(n1535), .OUT(n5343) );
  NAND2 U3465 ( .A(n5343), .B(n1534), .OUT(n4315) );
  NAND2 U3466 ( .A(n3118), .B(n4315), .OUT(n1637) );
  NAND2 U3467 ( .A(\mult_49/ab[17][10] ), .B(n1535), .OUT(n1636) );
  INV U3468 ( .IN(n1635), .OUT(n5344) );
  NAND2 U3469 ( .A(n5344), .B(n1634), .OUT(n4364) );
  NAND2 U3470 ( .A(n3193), .B(n4364), .OUT(n1741) );
  NAND2 U3471 ( .A(\mult_49/ab[18][10] ), .B(n1635), .OUT(n1740) );
  INV U3472 ( .IN(n1739), .OUT(n5345) );
  NAND2 U3473 ( .A(n5345), .B(n1738), .OUT(n4415) );
  NAND2 U3474 ( .A(n3271), .B(n4415), .OUT(n1849) );
  NAND2 U3475 ( .A(\mult_49/ab[19][10] ), .B(n1739), .OUT(n1848) );
  INV U3476 ( .IN(n1847), .OUT(n5346) );
  NAND2 U3477 ( .A(n5346), .B(n1846), .OUT(n4485) );
  NAND2 U3478 ( .A(n3352), .B(n4485), .OUT(n4841) );
  NAND2 U3479 ( .A(\mult_49/ab[20][10] ), .B(n1847), .OUT(n4486) );
  NAND2 U3480 ( .A(n5089), .B(n294), .OUT(n5347) );
  NAND2 U3481 ( .A(n2180), .B(n5347), .OUT(n521) );
  NAND2 U3482 ( .A(\mult_49/ab[2][9] ), .B(n291), .OUT(n520) );
  INV U3483 ( .IN(n519), .OUT(n5348) );
  NAND2 U3484 ( .A(n5348), .B(n518), .OUT(n3822) );
  NAND2 U3485 ( .A(n2356), .B(n3822), .OUT(n561) );
  NAND2 U3486 ( .A(\mult_49/ab[3][9] ), .B(n519), .OUT(n560) );
  INV U3487 ( .IN(n559), .OUT(n5349) );
  NAND2 U3488 ( .A(n5349), .B(n558), .OUT(n3841) );
  NAND2 U3489 ( .A(n2386), .B(n3841), .OUT(n605) );
  NAND2 U3490 ( .A(\mult_49/ab[4][9] ), .B(n559), .OUT(n604) );
  INV U3491 ( .IN(n603), .OUT(n5350) );
  NAND2 U3492 ( .A(n5350), .B(n602), .OUT(n3862) );
  NAND2 U3493 ( .A(n2419), .B(n3862), .OUT(n653) );
  NAND2 U3494 ( .A(\mult_49/ab[5][9] ), .B(n603), .OUT(n652) );
  INV U3495 ( .IN(n651), .OUT(n5351) );
  NAND2 U3496 ( .A(n5351), .B(n650), .OUT(n3885) );
  NAND2 U3497 ( .A(n2455), .B(n3885), .OUT(n705) );
  NAND2 U3498 ( .A(\mult_49/ab[6][9] ), .B(n651), .OUT(n704) );
  INV U3499 ( .IN(n703), .OUT(n5352) );
  NAND2 U3500 ( .A(n5352), .B(n702), .OUT(n3910) );
  NAND2 U3501 ( .A(n2494), .B(n3910), .OUT(n761) );
  NAND2 U3502 ( .A(\mult_49/ab[7][9] ), .B(n703), .OUT(n760) );
  INV U3503 ( .IN(n759), .OUT(n5353) );
  NAND2 U3504 ( .A(n5353), .B(n758), .OUT(n3937) );
  NAND2 U3505 ( .A(n2536), .B(n3937), .OUT(n821) );
  NAND2 U3506 ( .A(\mult_49/ab[8][9] ), .B(n759), .OUT(n820) );
  INV U3507 ( .IN(n819), .OUT(n5354) );
  NAND2 U3508 ( .A(n5354), .B(n818), .OUT(n3966) );
  NAND2 U3509 ( .A(n2581), .B(n3966), .OUT(n885) );
  NAND2 U3510 ( .A(\mult_49/ab[9][9] ), .B(n819), .OUT(n884) );
  INV U3511 ( .IN(n883), .OUT(n5355) );
  NAND2 U3512 ( .A(n5355), .B(n882), .OUT(n3997) );
  NAND2 U3513 ( .A(n2629), .B(n3997), .OUT(n953) );
  NAND2 U3514 ( .A(\mult_49/ab[10][9] ), .B(n883), .OUT(n952) );
  INV U3515 ( .IN(n951), .OUT(n5356) );
  NAND2 U3516 ( .A(n5356), .B(n950), .OUT(n4030) );
  NAND2 U3517 ( .A(n2680), .B(n4030), .OUT(n1025) );
  NAND2 U3518 ( .A(\mult_49/ab[11][9] ), .B(n951), .OUT(n1024) );
  INV U3519 ( .IN(n1023), .OUT(n5357) );
  NAND2 U3520 ( .A(n5357), .B(n1022), .OUT(n4065) );
  NAND2 U3521 ( .A(n2734), .B(n4065), .OUT(n1101) );
  NAND2 U3522 ( .A(\mult_49/ab[12][9] ), .B(n1023), .OUT(n1100) );
  INV U3523 ( .IN(n1099), .OUT(n5358) );
  NAND2 U3524 ( .A(n5358), .B(n1098), .OUT(n4102) );
  NAND2 U3525 ( .A(n2791), .B(n4102), .OUT(n1181) );
  NAND2 U3526 ( .A(\mult_49/ab[13][9] ), .B(n1099), .OUT(n1180) );
  INV U3527 ( .IN(n1179), .OUT(n5359) );
  NAND2 U3528 ( .A(n5359), .B(n1178), .OUT(n4141) );
  NAND2 U3529 ( .A(n2851), .B(n4141), .OUT(n1265) );
  NAND2 U3530 ( .A(\mult_49/ab[14][9] ), .B(n1179), .OUT(n1264) );
  INV U3531 ( .IN(n1263), .OUT(n5360) );
  NAND2 U3532 ( .A(n5360), .B(n1262), .OUT(n4182) );
  NAND2 U3533 ( .A(n2914), .B(n4182), .OUT(n1353) );
  NAND2 U3534 ( .A(\mult_49/ab[15][9] ), .B(n1263), .OUT(n1352) );
  INV U3535 ( .IN(n1351), .OUT(n5361) );
  NAND2 U3536 ( .A(n5361), .B(n1350), .OUT(n4225) );
  NAND2 U3537 ( .A(n2980), .B(n4225), .OUT(n1445) );
  NAND2 U3538 ( .A(\mult_49/ab[16][9] ), .B(n1351), .OUT(n1444) );
  INV U3539 ( .IN(n1443), .OUT(n5362) );
  NAND2 U3540 ( .A(n5362), .B(n1442), .OUT(n4270) );
  NAND2 U3541 ( .A(n3049), .B(n4270), .OUT(n1541) );
  NAND2 U3542 ( .A(\mult_49/ab[17][9] ), .B(n1443), .OUT(n1540) );
  INV U3543 ( .IN(n1539), .OUT(n5363) );
  NAND2 U3544 ( .A(n5363), .B(n1538), .OUT(n4317) );
  NAND2 U3545 ( .A(n3121), .B(n4317), .OUT(n1641) );
  NAND2 U3546 ( .A(\mult_49/ab[18][9] ), .B(n1539), .OUT(n1640) );
  INV U3547 ( .IN(n1639), .OUT(n5364) );
  NAND2 U3548 ( .A(n5364), .B(n1638), .OUT(n4366) );
  NAND2 U3549 ( .A(n3196), .B(n4366), .OUT(n1745) );
  NAND2 U3550 ( .A(\mult_49/ab[19][9] ), .B(n1639), .OUT(n1744) );
  INV U3551 ( .IN(n1743), .OUT(n5365) );
  NAND2 U3552 ( .A(n5365), .B(n1742), .OUT(n4417) );
  NAND2 U3553 ( .A(n3274), .B(n4417), .OUT(n1853) );
  NAND2 U3554 ( .A(\mult_49/ab[20][9] ), .B(n1743), .OUT(n1852) );
  INV U3555 ( .IN(n1851), .OUT(n5366) );
  NAND2 U3556 ( .A(n5366), .B(n1850), .OUT(n4488) );
  NAND2 U3557 ( .A(n3355), .B(n4488), .OUT(n4795) );
  NAND2 U3558 ( .A(\mult_49/ab[21][9] ), .B(n1851), .OUT(n4489) );
  NAND2 U3559 ( .A(n5100), .B(n299), .OUT(n3787) );
  NAND2 U3560 ( .A(n2183), .B(n3787), .OUT(n525) );
  NAND2 U3561 ( .A(\mult_49/ab[3][8] ), .B(n300), .OUT(n524) );
  INV U3562 ( .IN(n523), .OUT(n5367) );
  NAND2 U3563 ( .A(n5367), .B(n522), .OUT(n3824) );
  NAND2 U3564 ( .A(n2359), .B(n3824), .OUT(n565) );
  NAND2 U3565 ( .A(\mult_49/ab[4][8] ), .B(n523), .OUT(n564) );
  INV U3566 ( .IN(n563), .OUT(n5368) );
  NAND2 U3567 ( .A(n5368), .B(n562), .OUT(n3843) );
  NAND2 U3568 ( .A(n2389), .B(n3843), .OUT(n609) );
  NAND2 U3569 ( .A(\mult_49/ab[5][8] ), .B(n563), .OUT(n608) );
  INV U3570 ( .IN(n607), .OUT(n5369) );
  NAND2 U3571 ( .A(n5369), .B(n606), .OUT(n3864) );
  NAND2 U3572 ( .A(n2422), .B(n3864), .OUT(n657) );
  NAND2 U3573 ( .A(\mult_49/ab[6][8] ), .B(n607), .OUT(n656) );
  INV U3574 ( .IN(n655), .OUT(n5370) );
  NAND2 U3575 ( .A(n5370), .B(n654), .OUT(n3887) );
  NAND2 U3576 ( .A(n2458), .B(n3887), .OUT(n709) );
  NAND2 U3577 ( .A(\mult_49/ab[7][8] ), .B(n655), .OUT(n708) );
  INV U3578 ( .IN(n707), .OUT(n5371) );
  NAND2 U3579 ( .A(n5371), .B(n706), .OUT(n3912) );
  NAND2 U3580 ( .A(n2497), .B(n3912), .OUT(n765) );
  NAND2 U3581 ( .A(\mult_49/ab[8][8] ), .B(n707), .OUT(n764) );
  INV U3582 ( .IN(n763), .OUT(n5372) );
  NAND2 U3583 ( .A(n5372), .B(n762), .OUT(n3939) );
  NAND2 U3584 ( .A(n2539), .B(n3939), .OUT(n825) );
  NAND2 U3585 ( .A(\mult_49/ab[9][8] ), .B(n763), .OUT(n824) );
  INV U3586 ( .IN(n823), .OUT(n5373) );
  NAND2 U3587 ( .A(n5373), .B(n822), .OUT(n3968) );
  NAND2 U3588 ( .A(n2584), .B(n3968), .OUT(n889) );
  NAND2 U3589 ( .A(\mult_49/ab[10][8] ), .B(n823), .OUT(n888) );
  INV U3590 ( .IN(n887), .OUT(n5374) );
  NAND2 U3591 ( .A(n5374), .B(n886), .OUT(n3999) );
  NAND2 U3592 ( .A(n2632), .B(n3999), .OUT(n957) );
  NAND2 U3593 ( .A(\mult_49/ab[11][8] ), .B(n887), .OUT(n956) );
  INV U3594 ( .IN(n955), .OUT(n5375) );
  NAND2 U3595 ( .A(n5375), .B(n954), .OUT(n4032) );
  NAND2 U3596 ( .A(n2683), .B(n4032), .OUT(n1029) );
  NAND2 U3597 ( .A(\mult_49/ab[12][8] ), .B(n955), .OUT(n1028) );
  INV U3598 ( .IN(n1027), .OUT(n5376) );
  NAND2 U3599 ( .A(n5376), .B(n1026), .OUT(n4067) );
  NAND2 U3600 ( .A(n2737), .B(n4067), .OUT(n1105) );
  NAND2 U3601 ( .A(\mult_49/ab[13][8] ), .B(n1027), .OUT(n1104) );
  INV U3602 ( .IN(n1103), .OUT(n5377) );
  NAND2 U3603 ( .A(n5377), .B(n1102), .OUT(n4104) );
  NAND2 U3604 ( .A(n2794), .B(n4104), .OUT(n1185) );
  NAND2 U3605 ( .A(\mult_49/ab[14][8] ), .B(n1103), .OUT(n1184) );
  INV U3606 ( .IN(n1183), .OUT(n5378) );
  NAND2 U3607 ( .A(n5378), .B(n1182), .OUT(n4143) );
  NAND2 U3608 ( .A(n2854), .B(n4143), .OUT(n1269) );
  NAND2 U3609 ( .A(\mult_49/ab[15][8] ), .B(n1183), .OUT(n1268) );
  INV U3610 ( .IN(n1267), .OUT(n5379) );
  NAND2 U3611 ( .A(n5379), .B(n1266), .OUT(n4184) );
  NAND2 U3612 ( .A(n2917), .B(n4184), .OUT(n1357) );
  NAND2 U3613 ( .A(\mult_49/ab[16][8] ), .B(n1267), .OUT(n1356) );
  INV U3614 ( .IN(n1355), .OUT(n5380) );
  NAND2 U3615 ( .A(n5380), .B(n1354), .OUT(n4227) );
  NAND2 U3616 ( .A(n2983), .B(n4227), .OUT(n1449) );
  NAND2 U3617 ( .A(\mult_49/ab[17][8] ), .B(n1355), .OUT(n1448) );
  INV U3618 ( .IN(n1447), .OUT(n5381) );
  NAND2 U3619 ( .A(n5381), .B(n1446), .OUT(n4272) );
  NAND2 U3620 ( .A(n3052), .B(n4272), .OUT(n1545) );
  NAND2 U3621 ( .A(\mult_49/ab[18][8] ), .B(n1447), .OUT(n1544) );
  INV U3622 ( .IN(n1543), .OUT(n5382) );
  NAND2 U3623 ( .A(n5382), .B(n1542), .OUT(n4319) );
  NAND2 U3624 ( .A(n3124), .B(n4319), .OUT(n1645) );
  NAND2 U3625 ( .A(\mult_49/ab[19][8] ), .B(n1543), .OUT(n1644) );
  INV U3626 ( .IN(n1643), .OUT(n5383) );
  NAND2 U3627 ( .A(n5383), .B(n1642), .OUT(n4368) );
  NAND2 U3628 ( .A(n3199), .B(n4368), .OUT(n1749) );
  NAND2 U3629 ( .A(\mult_49/ab[20][8] ), .B(n1643), .OUT(n1748) );
  INV U3630 ( .IN(n1747), .OUT(n5384) );
  NAND2 U3631 ( .A(n5384), .B(n1746), .OUT(n4419) );
  NAND2 U3632 ( .A(n3277), .B(n4419), .OUT(n1857) );
  NAND2 U3633 ( .A(\mult_49/ab[21][8] ), .B(n1747), .OUT(n1856) );
  INV U3634 ( .IN(n1855), .OUT(n5385) );
  NAND2 U3635 ( .A(n5385), .B(n1854), .OUT(n4491) );
  NAND2 U3636 ( .A(n3358), .B(n4491), .OUT(n4797) );
  NAND2 U3637 ( .A(\mult_49/ab[22][8] ), .B(n1855), .OUT(n4492) );
  NAND2 U3638 ( .A(n5103), .B(n311), .OUT(n3789) );
  NAND2 U3639 ( .A(n2189), .B(n3789), .OUT(n529) );
  NAND2 U3640 ( .A(\mult_49/ab[4][7] ), .B(n312), .OUT(n528) );
  INV U3641 ( .IN(n527), .OUT(n5386) );
  NAND2 U3642 ( .A(n5386), .B(n526), .OUT(n3826) );
  NAND2 U3643 ( .A(n2362), .B(n3826), .OUT(n569) );
  NAND2 U3644 ( .A(\mult_49/ab[5][7] ), .B(n527), .OUT(n568) );
  INV U3645 ( .IN(n567), .OUT(n5387) );
  NAND2 U3646 ( .A(n5387), .B(n566), .OUT(n3845) );
  NAND2 U3647 ( .A(n2392), .B(n3845), .OUT(n613) );
  NAND2 U3648 ( .A(\mult_49/ab[6][7] ), .B(n567), .OUT(n612) );
  INV U3649 ( .IN(n611), .OUT(n5388) );
  NAND2 U3650 ( .A(n5388), .B(n610), .OUT(n3866) );
  NAND2 U3651 ( .A(n2425), .B(n3866), .OUT(n661) );
  NAND2 U3652 ( .A(\mult_49/ab[7][7] ), .B(n611), .OUT(n660) );
  INV U3653 ( .IN(n659), .OUT(n5389) );
  NAND2 U3654 ( .A(n5389), .B(n658), .OUT(n3889) );
  NAND2 U3655 ( .A(n2461), .B(n3889), .OUT(n713) );
  NAND2 U3656 ( .A(\mult_49/ab[8][7] ), .B(n659), .OUT(n712) );
  INV U3657 ( .IN(n711), .OUT(n5390) );
  NAND2 U3658 ( .A(n5390), .B(n710), .OUT(n3914) );
  NAND2 U3659 ( .A(n2500), .B(n3914), .OUT(n769) );
  NAND2 U3660 ( .A(\mult_49/ab[9][7] ), .B(n711), .OUT(n768) );
  INV U3661 ( .IN(n767), .OUT(n5391) );
  NAND2 U3662 ( .A(n5391), .B(n766), .OUT(n3941) );
  NAND2 U3663 ( .A(n2542), .B(n3941), .OUT(n829) );
  NAND2 U3664 ( .A(\mult_49/ab[10][7] ), .B(n767), .OUT(n828) );
  INV U3665 ( .IN(n827), .OUT(n5392) );
  NAND2 U3666 ( .A(n5392), .B(n826), .OUT(n3970) );
  NAND2 U3667 ( .A(n2587), .B(n3970), .OUT(n893) );
  NAND2 U3668 ( .A(\mult_49/ab[11][7] ), .B(n827), .OUT(n892) );
  INV U3669 ( .IN(n891), .OUT(n5393) );
  NAND2 U3670 ( .A(n5393), .B(n890), .OUT(n4001) );
  NAND2 U3671 ( .A(n2635), .B(n4001), .OUT(n961) );
  NAND2 U3672 ( .A(\mult_49/ab[12][7] ), .B(n891), .OUT(n960) );
  INV U3673 ( .IN(n959), .OUT(n5394) );
  NAND2 U3674 ( .A(n5394), .B(n958), .OUT(n4034) );
  NAND2 U3675 ( .A(n2686), .B(n4034), .OUT(n1033) );
  NAND2 U3676 ( .A(\mult_49/ab[13][7] ), .B(n959), .OUT(n1032) );
  INV U3677 ( .IN(n1031), .OUT(n5395) );
  NAND2 U3678 ( .A(n5395), .B(n1030), .OUT(n4069) );
  NAND2 U3679 ( .A(n2740), .B(n4069), .OUT(n1109) );
  NAND2 U3680 ( .A(\mult_49/ab[14][7] ), .B(n1031), .OUT(n1108) );
  INV U3681 ( .IN(n1107), .OUT(n5396) );
  NAND2 U3682 ( .A(n5396), .B(n1106), .OUT(n4106) );
  NAND2 U3683 ( .A(n2797), .B(n4106), .OUT(n1189) );
  NAND2 U3684 ( .A(\mult_49/ab[15][7] ), .B(n1107), .OUT(n1188) );
  INV U3685 ( .IN(n1187), .OUT(n5397) );
  NAND2 U3686 ( .A(n5397), .B(n1186), .OUT(n4145) );
  NAND2 U3687 ( .A(n2857), .B(n4145), .OUT(n1273) );
  NAND2 U3688 ( .A(\mult_49/ab[16][7] ), .B(n1187), .OUT(n1272) );
  INV U3689 ( .IN(n1271), .OUT(n5398) );
  NAND2 U3690 ( .A(n5398), .B(n1270), .OUT(n4186) );
  NAND2 U3691 ( .A(n2920), .B(n4186), .OUT(n1361) );
  NAND2 U3692 ( .A(\mult_49/ab[17][7] ), .B(n1271), .OUT(n1360) );
  INV U3693 ( .IN(n1359), .OUT(n5399) );
  NAND2 U3694 ( .A(n5399), .B(n1358), .OUT(n4229) );
  NAND2 U3695 ( .A(n2986), .B(n4229), .OUT(n1453) );
  NAND2 U3696 ( .A(\mult_49/ab[18][7] ), .B(n1359), .OUT(n1452) );
  INV U3697 ( .IN(n1451), .OUT(n5400) );
  NAND2 U3698 ( .A(n5400), .B(n1450), .OUT(n4274) );
  NAND2 U3699 ( .A(n3055), .B(n4274), .OUT(n1549) );
  NAND2 U3700 ( .A(\mult_49/ab[19][7] ), .B(n1451), .OUT(n1548) );
  INV U3701 ( .IN(n1547), .OUT(n5401) );
  NAND2 U3702 ( .A(n5401), .B(n1546), .OUT(n4321) );
  NAND2 U3703 ( .A(n3127), .B(n4321), .OUT(n1649) );
  NAND2 U3704 ( .A(\mult_49/ab[20][7] ), .B(n1547), .OUT(n1648) );
  INV U3705 ( .IN(n1647), .OUT(n5402) );
  NAND2 U3706 ( .A(n5402), .B(n1646), .OUT(n4370) );
  NAND2 U3707 ( .A(n3202), .B(n4370), .OUT(n1753) );
  NAND2 U3708 ( .A(\mult_49/ab[21][7] ), .B(n1647), .OUT(n1752) );
  INV U3709 ( .IN(n1751), .OUT(n5403) );
  NAND2 U3710 ( .A(n5403), .B(n1750), .OUT(n4421) );
  NAND2 U3711 ( .A(n3280), .B(n4421), .OUT(n1861) );
  NAND2 U3712 ( .A(\mult_49/ab[22][7] ), .B(n1751), .OUT(n1860) );
  INV U3713 ( .IN(n1859), .OUT(n5404) );
  NAND2 U3714 ( .A(n5404), .B(n1858), .OUT(n4494) );
  NAND2 U3715 ( .A(n3361), .B(n4494), .OUT(n4801) );
  NAND2 U3716 ( .A(\mult_49/ab[23][7] ), .B(n1859), .OUT(n4495) );
  NAND2 U3717 ( .A(n5107), .B(n327), .OUT(n3791) );
  NAND2 U3718 ( .A(n2198), .B(n3791), .OUT(n533) );
  NAND2 U3719 ( .A(\mult_49/ab[5][6] ), .B(n328), .OUT(n532) );
  INV U3720 ( .IN(n531), .OUT(n5405) );
  NAND2 U3721 ( .A(n5405), .B(n530), .OUT(n3828) );
  NAND2 U3722 ( .A(n2365), .B(n3828), .OUT(n573) );
  NAND2 U3723 ( .A(\mult_49/ab[6][6] ), .B(n531), .OUT(n572) );
  INV U3724 ( .IN(n571), .OUT(n5406) );
  NAND2 U3725 ( .A(n5406), .B(n570), .OUT(n3847) );
  NAND2 U3726 ( .A(n2395), .B(n3847), .OUT(n617) );
  NAND2 U3727 ( .A(\mult_49/ab[7][6] ), .B(n571), .OUT(n616) );
  INV U3728 ( .IN(n615), .OUT(n5407) );
  NAND2 U3729 ( .A(n5407), .B(n614), .OUT(n3868) );
  NAND2 U3730 ( .A(n2428), .B(n3868), .OUT(n665) );
  NAND2 U3731 ( .A(\mult_49/ab[8][6] ), .B(n615), .OUT(n664) );
  INV U3732 ( .IN(n663), .OUT(n5408) );
  NAND2 U3733 ( .A(n5408), .B(n662), .OUT(n3891) );
  NAND2 U3734 ( .A(n2464), .B(n3891), .OUT(n717) );
  NAND2 U3735 ( .A(\mult_49/ab[9][6] ), .B(n663), .OUT(n716) );
  INV U3736 ( .IN(n715), .OUT(n5409) );
  NAND2 U3737 ( .A(n5409), .B(n714), .OUT(n3916) );
  NAND2 U3738 ( .A(n2503), .B(n3916), .OUT(n773) );
  NAND2 U3739 ( .A(\mult_49/ab[10][6] ), .B(n715), .OUT(n772) );
  INV U3740 ( .IN(n771), .OUT(n5410) );
  NAND2 U3741 ( .A(n5410), .B(n770), .OUT(n3943) );
  NAND2 U3742 ( .A(n2545), .B(n3943), .OUT(n833) );
  NAND2 U3743 ( .A(\mult_49/ab[11][6] ), .B(n771), .OUT(n832) );
  INV U3744 ( .IN(n831), .OUT(n5411) );
  NAND2 U3745 ( .A(n5411), .B(n830), .OUT(n3972) );
  NAND2 U3746 ( .A(n2590), .B(n3972), .OUT(n897) );
  NAND2 U3747 ( .A(\mult_49/ab[12][6] ), .B(n831), .OUT(n896) );
  INV U3748 ( .IN(n895), .OUT(n5412) );
  NAND2 U3749 ( .A(n5412), .B(n894), .OUT(n4003) );
  NAND2 U3750 ( .A(n2638), .B(n4003), .OUT(n965) );
  NAND2 U3751 ( .A(\mult_49/ab[13][6] ), .B(n895), .OUT(n964) );
  INV U3752 ( .IN(n963), .OUT(n5413) );
  NAND2 U3753 ( .A(n5413), .B(n962), .OUT(n4036) );
  NAND2 U3754 ( .A(n2689), .B(n4036), .OUT(n1037) );
  NAND2 U3755 ( .A(\mult_49/ab[14][6] ), .B(n963), .OUT(n1036) );
  INV U3756 ( .IN(n1035), .OUT(n5414) );
  NAND2 U3757 ( .A(n5414), .B(n1034), .OUT(n4071) );
  NAND2 U3758 ( .A(n2743), .B(n4071), .OUT(n1113) );
  NAND2 U3759 ( .A(\mult_49/ab[15][6] ), .B(n1035), .OUT(n1112) );
  INV U3760 ( .IN(n1111), .OUT(n5415) );
  NAND2 U3761 ( .A(n5415), .B(n1110), .OUT(n4108) );
  NAND2 U3762 ( .A(n2800), .B(n4108), .OUT(n1193) );
  NAND2 U3763 ( .A(\mult_49/ab[16][6] ), .B(n1111), .OUT(n1192) );
  INV U3764 ( .IN(n1191), .OUT(n5416) );
  NAND2 U3765 ( .A(n5416), .B(n1190), .OUT(n4147) );
  NAND2 U3766 ( .A(n2860), .B(n4147), .OUT(n1277) );
  NAND2 U3767 ( .A(\mult_49/ab[17][6] ), .B(n1191), .OUT(n1276) );
  INV U3768 ( .IN(n1275), .OUT(n5417) );
  NAND2 U3769 ( .A(n5417), .B(n1274), .OUT(n4188) );
  NAND2 U3770 ( .A(n2923), .B(n4188), .OUT(n1365) );
  NAND2 U3771 ( .A(\mult_49/ab[18][6] ), .B(n1275), .OUT(n1364) );
  INV U3772 ( .IN(n1363), .OUT(n5418) );
  NAND2 U3773 ( .A(n5418), .B(n1362), .OUT(n4231) );
  NAND2 U3774 ( .A(n2989), .B(n4231), .OUT(n1457) );
  NAND2 U3775 ( .A(\mult_49/ab[19][6] ), .B(n1363), .OUT(n1456) );
  INV U3776 ( .IN(n1455), .OUT(n5419) );
  NAND2 U3777 ( .A(n5419), .B(n1454), .OUT(n4276) );
  NAND2 U3778 ( .A(n3058), .B(n4276), .OUT(n1553) );
  NAND2 U3779 ( .A(\mult_49/ab[20][6] ), .B(n1455), .OUT(n1552) );
  INV U3780 ( .IN(n1551), .OUT(n5420) );
  NAND2 U3781 ( .A(n5420), .B(n1550), .OUT(n4323) );
  NAND2 U3782 ( .A(n3130), .B(n4323), .OUT(n1653) );
  NAND2 U3783 ( .A(\mult_49/ab[21][6] ), .B(n1551), .OUT(n1652) );
  INV U3784 ( .IN(n1651), .OUT(n5421) );
  NAND2 U3785 ( .A(n5421), .B(n1650), .OUT(n4372) );
  NAND2 U3786 ( .A(n3205), .B(n4372), .OUT(n1757) );
  NAND2 U3787 ( .A(\mult_49/ab[22][6] ), .B(n1651), .OUT(n1756) );
  INV U3788 ( .IN(n1755), .OUT(n5422) );
  NAND2 U3789 ( .A(n5422), .B(n1754), .OUT(n4423) );
  NAND2 U3790 ( .A(n3283), .B(n4423), .OUT(n1865) );
  NAND2 U3791 ( .A(\mult_49/ab[23][6] ), .B(n1755), .OUT(n1864) );
  INV U3792 ( .IN(n1863), .OUT(n5423) );
  NAND2 U3793 ( .A(n5423), .B(n1862), .OUT(n4497) );
  NAND2 U3794 ( .A(n3364), .B(n4497), .OUT(n4793) );
  NAND2 U3795 ( .A(\mult_49/ab[24][6] ), .B(n1863), .OUT(n4498) );
  NAND2 U3796 ( .A(n5112), .B(n347), .OUT(n3793) );
  NAND2 U3797 ( .A(n2210), .B(n3793), .OUT(n537) );
  NAND2 U3798 ( .A(\mult_49/ab[6][5] ), .B(n348), .OUT(n536) );
  INV U3799 ( .IN(n535), .OUT(n5424) );
  NAND2 U3800 ( .A(n5424), .B(n534), .OUT(n3830) );
  NAND2 U3801 ( .A(n2368), .B(n3830), .OUT(n577) );
  NAND2 U3802 ( .A(\mult_49/ab[7][5] ), .B(n535), .OUT(n576) );
  INV U3803 ( .IN(n575), .OUT(n5425) );
  NAND2 U3804 ( .A(n5425), .B(n574), .OUT(n3849) );
  NAND2 U3805 ( .A(n2398), .B(n3849), .OUT(n621) );
  NAND2 U3806 ( .A(\mult_49/ab[8][5] ), .B(n575), .OUT(n620) );
  INV U3807 ( .IN(n619), .OUT(n5426) );
  NAND2 U3808 ( .A(n5426), .B(n618), .OUT(n3870) );
  NAND2 U3809 ( .A(n2431), .B(n3870), .OUT(n669) );
  NAND2 U3810 ( .A(\mult_49/ab[9][5] ), .B(n619), .OUT(n668) );
  INV U3811 ( .IN(n667), .OUT(n5427) );
  NAND2 U3812 ( .A(n5427), .B(n666), .OUT(n3893) );
  NAND2 U3813 ( .A(n2467), .B(n3893), .OUT(n721) );
  NAND2 U3814 ( .A(\mult_49/ab[10][5] ), .B(n667), .OUT(n720) );
  INV U3815 ( .IN(n719), .OUT(n5428) );
  NAND2 U3816 ( .A(n5428), .B(n718), .OUT(n3918) );
  NAND2 U3817 ( .A(n2506), .B(n3918), .OUT(n777) );
  NAND2 U3818 ( .A(\mult_49/ab[11][5] ), .B(n719), .OUT(n776) );
  INV U3819 ( .IN(n775), .OUT(n5429) );
  NAND2 U3820 ( .A(n5429), .B(n774), .OUT(n3945) );
  NAND2 U3821 ( .A(n2548), .B(n3945), .OUT(n837) );
  NAND2 U3822 ( .A(\mult_49/ab[12][5] ), .B(n775), .OUT(n836) );
  INV U3823 ( .IN(n835), .OUT(n5430) );
  NAND2 U3824 ( .A(n5430), .B(n834), .OUT(n3974) );
  NAND2 U3825 ( .A(n2593), .B(n3974), .OUT(n901) );
  NAND2 U3826 ( .A(\mult_49/ab[13][5] ), .B(n835), .OUT(n900) );
  INV U3827 ( .IN(n899), .OUT(n5431) );
  NAND2 U3828 ( .A(n5431), .B(n898), .OUT(n4005) );
  NAND2 U3829 ( .A(n2641), .B(n4005), .OUT(n969) );
  NAND2 U3830 ( .A(\mult_49/ab[14][5] ), .B(n899), .OUT(n968) );
  INV U3831 ( .IN(n967), .OUT(n5432) );
  NAND2 U3832 ( .A(n5432), .B(n966), .OUT(n4038) );
  NAND2 U3833 ( .A(n2692), .B(n4038), .OUT(n1041) );
  NAND2 U3834 ( .A(\mult_49/ab[15][5] ), .B(n967), .OUT(n1040) );
  INV U3835 ( .IN(n1039), .OUT(n5433) );
  NAND2 U3836 ( .A(n5433), .B(n1038), .OUT(n4073) );
  NAND2 U3837 ( .A(n2746), .B(n4073), .OUT(n1117) );
  NAND2 U3838 ( .A(\mult_49/ab[16][5] ), .B(n1039), .OUT(n1116) );
  INV U3839 ( .IN(n1115), .OUT(n5434) );
  NAND2 U3840 ( .A(n5434), .B(n1114), .OUT(n4110) );
  NAND2 U3841 ( .A(n2803), .B(n4110), .OUT(n1197) );
  NAND2 U3842 ( .A(\mult_49/ab[17][5] ), .B(n1115), .OUT(n1196) );
  INV U3843 ( .IN(n1195), .OUT(n5435) );
  NAND2 U3844 ( .A(n5435), .B(n1194), .OUT(n4149) );
  NAND2 U3845 ( .A(n2863), .B(n4149), .OUT(n1281) );
  NAND2 U3846 ( .A(\mult_49/ab[18][5] ), .B(n1195), .OUT(n1280) );
  INV U3847 ( .IN(n1279), .OUT(n5436) );
  NAND2 U3848 ( .A(n5436), .B(n1278), .OUT(n4190) );
  NAND2 U3849 ( .A(n2926), .B(n4190), .OUT(n1369) );
  NAND2 U3850 ( .A(\mult_49/ab[19][5] ), .B(n1279), .OUT(n1368) );
  INV U3851 ( .IN(n1367), .OUT(n5437) );
  NAND2 U3852 ( .A(n5437), .B(n1366), .OUT(n4233) );
  NAND2 U3853 ( .A(n2992), .B(n4233), .OUT(n1461) );
  NAND2 U3854 ( .A(\mult_49/ab[20][5] ), .B(n1367), .OUT(n1460) );
  INV U3855 ( .IN(n1459), .OUT(n5438) );
  NAND2 U3856 ( .A(n5438), .B(n1458), .OUT(n4278) );
  NAND2 U3857 ( .A(n3061), .B(n4278), .OUT(n1557) );
  NAND2 U3858 ( .A(\mult_49/ab[21][5] ), .B(n1459), .OUT(n1556) );
  INV U3859 ( .IN(n1555), .OUT(n5439) );
  NAND2 U3860 ( .A(n5439), .B(n1554), .OUT(n4325) );
  NAND2 U3861 ( .A(n3133), .B(n4325), .OUT(n1657) );
  NAND2 U3862 ( .A(\mult_49/ab[22][5] ), .B(n1555), .OUT(n1656) );
  INV U3863 ( .IN(n1655), .OUT(n5440) );
  NAND2 U3864 ( .A(n5440), .B(n1654), .OUT(n4374) );
  NAND2 U3865 ( .A(n3208), .B(n4374), .OUT(n1761) );
  NAND2 U3866 ( .A(\mult_49/ab[23][5] ), .B(n1655), .OUT(n1760) );
  INV U3867 ( .IN(n1759), .OUT(n5441) );
  NAND2 U3868 ( .A(n5441), .B(n1758), .OUT(n4425) );
  NAND2 U3869 ( .A(n3286), .B(n4425), .OUT(n1869) );
  NAND2 U3870 ( .A(\mult_49/ab[24][5] ), .B(n1759), .OUT(n1868) );
  INV U3871 ( .IN(n1867), .OUT(n5442) );
  NAND2 U3872 ( .A(n5442), .B(n1866), .OUT(n4500) );
  NAND2 U3873 ( .A(n3367), .B(n4500), .OUT(n4843) );
  NAND2 U3874 ( .A(\mult_49/ab[25][5] ), .B(n1867), .OUT(n4501) );
  NAND2 U3875 ( .A(n5118), .B(n371), .OUT(n3795) );
  NAND2 U3876 ( .A(n2225), .B(n3795), .OUT(n541) );
  NAND2 U3877 ( .A(\mult_49/ab[7][4] ), .B(n372), .OUT(n540) );
  INV U3878 ( .IN(n539), .OUT(n5443) );
  NAND2 U3879 ( .A(n5443), .B(n538), .OUT(n3832) );
  NAND2 U3880 ( .A(n2371), .B(n3832), .OUT(n581) );
  NAND2 U3881 ( .A(\mult_49/ab[8][4] ), .B(n539), .OUT(n580) );
  INV U3882 ( .IN(n579), .OUT(n5444) );
  NAND2 U3883 ( .A(n5444), .B(n578), .OUT(n3851) );
  NAND2 U3884 ( .A(n2401), .B(n3851), .OUT(n625) );
  NAND2 U3885 ( .A(\mult_49/ab[9][4] ), .B(n579), .OUT(n624) );
  INV U3886 ( .IN(n623), .OUT(n5445) );
  NAND2 U3887 ( .A(n5445), .B(n622), .OUT(n3872) );
  NAND2 U3888 ( .A(n2434), .B(n3872), .OUT(n673) );
  NAND2 U3889 ( .A(\mult_49/ab[10][4] ), .B(n623), .OUT(n672) );
  INV U3890 ( .IN(n671), .OUT(n5446) );
  NAND2 U3891 ( .A(n5446), .B(n670), .OUT(n3895) );
  NAND2 U3892 ( .A(n2470), .B(n3895), .OUT(n725) );
  NAND2 U3893 ( .A(\mult_49/ab[11][4] ), .B(n671), .OUT(n724) );
  INV U3894 ( .IN(n723), .OUT(n5447) );
  NAND2 U3895 ( .A(n5447), .B(n722), .OUT(n3920) );
  NAND2 U3896 ( .A(n2509), .B(n3920), .OUT(n781) );
  NAND2 U3897 ( .A(\mult_49/ab[12][4] ), .B(n723), .OUT(n780) );
  INV U3898 ( .IN(n779), .OUT(n5448) );
  NAND2 U3899 ( .A(n5448), .B(n778), .OUT(n3947) );
  NAND2 U3900 ( .A(n2551), .B(n3947), .OUT(n841) );
  NAND2 U3901 ( .A(\mult_49/ab[13][4] ), .B(n779), .OUT(n840) );
  INV U3902 ( .IN(n839), .OUT(n5449) );
  NAND2 U3903 ( .A(n5449), .B(n838), .OUT(n3976) );
  NAND2 U3904 ( .A(n2596), .B(n3976), .OUT(n905) );
  NAND2 U3905 ( .A(\mult_49/ab[14][4] ), .B(n839), .OUT(n904) );
  INV U3906 ( .IN(n903), .OUT(n5450) );
  NAND2 U3907 ( .A(n5450), .B(n902), .OUT(n4007) );
  NAND2 U3908 ( .A(n2644), .B(n4007), .OUT(n973) );
  NAND2 U3909 ( .A(\mult_49/ab[15][4] ), .B(n903), .OUT(n972) );
  INV U3910 ( .IN(n971), .OUT(n5451) );
  NAND2 U3911 ( .A(n5451), .B(n970), .OUT(n4040) );
  NAND2 U3912 ( .A(n2695), .B(n4040), .OUT(n1045) );
  NAND2 U3913 ( .A(\mult_49/ab[16][4] ), .B(n971), .OUT(n1044) );
  INV U3914 ( .IN(n1043), .OUT(n5452) );
  NAND2 U3915 ( .A(n5452), .B(n1042), .OUT(n4075) );
  NAND2 U3916 ( .A(n2749), .B(n4075), .OUT(n1121) );
  NAND2 U3917 ( .A(\mult_49/ab[17][4] ), .B(n1043), .OUT(n1120) );
  INV U3918 ( .IN(n1119), .OUT(n5453) );
  NAND2 U3919 ( .A(n5453), .B(n1118), .OUT(n4112) );
  NAND2 U3920 ( .A(n2806), .B(n4112), .OUT(n1201) );
  NAND2 U3921 ( .A(\mult_49/ab[18][4] ), .B(n1119), .OUT(n1200) );
  INV U3922 ( .IN(n1199), .OUT(n5454) );
  NAND2 U3923 ( .A(n5454), .B(n1198), .OUT(n4151) );
  NAND2 U3924 ( .A(n2866), .B(n4151), .OUT(n1285) );
  NAND2 U3925 ( .A(\mult_49/ab[19][4] ), .B(n1199), .OUT(n1284) );
  INV U3926 ( .IN(n1283), .OUT(n5455) );
  NAND2 U3927 ( .A(n5455), .B(n1282), .OUT(n4192) );
  NAND2 U3928 ( .A(n2929), .B(n4192), .OUT(n1373) );
  NAND2 U3929 ( .A(\mult_49/ab[20][4] ), .B(n1283), .OUT(n1372) );
  INV U3930 ( .IN(n1371), .OUT(n5456) );
  NAND2 U3931 ( .A(n5456), .B(n1370), .OUT(n4235) );
  NAND2 U3932 ( .A(n2995), .B(n4235), .OUT(n1465) );
  NAND2 U3933 ( .A(\mult_49/ab[21][4] ), .B(n1371), .OUT(n1464) );
  INV U3934 ( .IN(n1463), .OUT(n5457) );
  NAND2 U3935 ( .A(n5457), .B(n1462), .OUT(n4280) );
  NAND2 U3936 ( .A(n3064), .B(n4280), .OUT(n1561) );
  NAND2 U3937 ( .A(\mult_49/ab[22][4] ), .B(n1463), .OUT(n1560) );
  INV U3938 ( .IN(n1559), .OUT(n5458) );
  NAND2 U3939 ( .A(n5458), .B(n1558), .OUT(n4327) );
  NAND2 U3940 ( .A(n3136), .B(n4327), .OUT(n1661) );
  NAND2 U3941 ( .A(\mult_49/ab[23][4] ), .B(n1559), .OUT(n1660) );
  INV U3942 ( .IN(n1659), .OUT(n5459) );
  NAND2 U3943 ( .A(n5459), .B(n1658), .OUT(n4376) );
  NAND2 U3944 ( .A(n3211), .B(n4376), .OUT(n1765) );
  NAND2 U3945 ( .A(\mult_49/ab[24][4] ), .B(n1659), .OUT(n1764) );
  INV U3946 ( .IN(n1763), .OUT(n5460) );
  NAND2 U3947 ( .A(n5460), .B(n1762), .OUT(n4427) );
  NAND2 U3948 ( .A(n3289), .B(n4427), .OUT(n1873) );
  NAND2 U3949 ( .A(\mult_49/ab[25][4] ), .B(n1763), .OUT(n1872) );
  INV U3950 ( .IN(n1871), .OUT(n5461) );
  NAND2 U3951 ( .A(n5461), .B(n1870), .OUT(n4503) );
  NAND2 U3952 ( .A(n3370), .B(n4503), .OUT(n4845) );
  NAND2 U3953 ( .A(\mult_49/ab[26][4] ), .B(n1871), .OUT(n4504) );
  NAND2 U3954 ( .A(n5125), .B(n399), .OUT(n3797) );
  NAND2 U3955 ( .A(n2243), .B(n3797), .OUT(n545) );
  NAND2 U3956 ( .A(\mult_49/ab[8][3] ), .B(n400), .OUT(n544) );
  INV U3957 ( .IN(n543), .OUT(n5462) );
  NAND2 U3958 ( .A(n5462), .B(n542), .OUT(n3834) );
  NAND2 U3959 ( .A(n2374), .B(n3834), .OUT(n585) );
  NAND2 U3960 ( .A(\mult_49/ab[9][3] ), .B(n543), .OUT(n584) );
  INV U3961 ( .IN(n583), .OUT(n5463) );
  NAND2 U3962 ( .A(n5463), .B(n582), .OUT(n3853) );
  NAND2 U3963 ( .A(n2404), .B(n3853), .OUT(n629) );
  NAND2 U3964 ( .A(\mult_49/ab[10][3] ), .B(n583), .OUT(n628) );
  INV U3965 ( .IN(n627), .OUT(n5464) );
  NAND2 U3966 ( .A(n5464), .B(n626), .OUT(n3874) );
  NAND2 U3967 ( .A(n2437), .B(n3874), .OUT(n677) );
  NAND2 U3968 ( .A(\mult_49/ab[11][3] ), .B(n627), .OUT(n676) );
  INV U3969 ( .IN(n675), .OUT(n5465) );
  NAND2 U3970 ( .A(n5465), .B(n674), .OUT(n3897) );
  NAND2 U3971 ( .A(n2473), .B(n3897), .OUT(n729) );
  NAND2 U3972 ( .A(\mult_49/ab[12][3] ), .B(n675), .OUT(n728) );
  INV U3973 ( .IN(n727), .OUT(n5466) );
  NAND2 U3974 ( .A(n5466), .B(n726), .OUT(n3922) );
  NAND2 U3975 ( .A(n2512), .B(n3922), .OUT(n785) );
  NAND2 U3976 ( .A(\mult_49/ab[13][3] ), .B(n727), .OUT(n784) );
  INV U3977 ( .IN(n783), .OUT(n5467) );
  NAND2 U3978 ( .A(n5467), .B(n782), .OUT(n3949) );
  NAND2 U3979 ( .A(n2554), .B(n3949), .OUT(n845) );
  NAND2 U3980 ( .A(\mult_49/ab[14][3] ), .B(n783), .OUT(n844) );
  INV U3981 ( .IN(n843), .OUT(n5468) );
  NAND2 U3982 ( .A(n5468), .B(n842), .OUT(n3978) );
  NAND2 U3983 ( .A(n2599), .B(n3978), .OUT(n909) );
  NAND2 U3984 ( .A(\mult_49/ab[15][3] ), .B(n843), .OUT(n908) );
  INV U3985 ( .IN(n907), .OUT(n5469) );
  NAND2 U3986 ( .A(n5469), .B(n906), .OUT(n4009) );
  NAND2 U3987 ( .A(n2647), .B(n4009), .OUT(n977) );
  NAND2 U3988 ( .A(\mult_49/ab[16][3] ), .B(n907), .OUT(n976) );
  INV U3989 ( .IN(n975), .OUT(n5470) );
  NAND2 U3990 ( .A(n5470), .B(n974), .OUT(n4042) );
  NAND2 U3991 ( .A(n2698), .B(n4042), .OUT(n1049) );
  NAND2 U3992 ( .A(\mult_49/ab[17][3] ), .B(n975), .OUT(n1048) );
  INV U3993 ( .IN(n1047), .OUT(n5471) );
  NAND2 U3994 ( .A(n5471), .B(n1046), .OUT(n4077) );
  NAND2 U3995 ( .A(n2752), .B(n4077), .OUT(n1125) );
  NAND2 U3996 ( .A(\mult_49/ab[18][3] ), .B(n1047), .OUT(n1124) );
  INV U3997 ( .IN(n1123), .OUT(n5472) );
  NAND2 U3998 ( .A(n5472), .B(n1122), .OUT(n4114) );
  NAND2 U3999 ( .A(n2809), .B(n4114), .OUT(n1205) );
  NAND2 U4000 ( .A(\mult_49/ab[19][3] ), .B(n1123), .OUT(n1204) );
  INV U4001 ( .IN(n1203), .OUT(n5473) );
  NAND2 U4002 ( .A(n5473), .B(n1202), .OUT(n4153) );
  NAND2 U4003 ( .A(n2869), .B(n4153), .OUT(n1289) );
  NAND2 U4004 ( .A(\mult_49/ab[20][3] ), .B(n1203), .OUT(n1288) );
  INV U4005 ( .IN(n1287), .OUT(n5474) );
  NAND2 U4006 ( .A(n5474), .B(n1286), .OUT(n4194) );
  NAND2 U4007 ( .A(n2932), .B(n4194), .OUT(n1377) );
  NAND2 U4008 ( .A(\mult_49/ab[21][3] ), .B(n1287), .OUT(n1376) );
  INV U4009 ( .IN(n1375), .OUT(n5475) );
  NAND2 U4010 ( .A(n5475), .B(n1374), .OUT(n4237) );
  NAND2 U4011 ( .A(n2998), .B(n4237), .OUT(n1469) );
  NAND2 U4012 ( .A(\mult_49/ab[22][3] ), .B(n1375), .OUT(n1468) );
  INV U4013 ( .IN(n1467), .OUT(n5476) );
  NAND2 U4014 ( .A(n5476), .B(n1466), .OUT(n4282) );
  NAND2 U4015 ( .A(n3067), .B(n4282), .OUT(n1565) );
  NAND2 U4016 ( .A(\mult_49/ab[23][3] ), .B(n1467), .OUT(n1564) );
  INV U4017 ( .IN(n1563), .OUT(n5477) );
  NAND2 U4018 ( .A(n5477), .B(n1562), .OUT(n4329) );
  NAND2 U4019 ( .A(n3139), .B(n4329), .OUT(n1665) );
  NAND2 U4020 ( .A(\mult_49/ab[24][3] ), .B(n1563), .OUT(n1664) );
  INV U4021 ( .IN(n1663), .OUT(n5478) );
  NAND2 U4022 ( .A(n5478), .B(n1662), .OUT(n4378) );
  NAND2 U4023 ( .A(n3214), .B(n4378), .OUT(n1769) );
  NAND2 U4024 ( .A(\mult_49/ab[25][3] ), .B(n1663), .OUT(n1768) );
  INV U4025 ( .IN(n1767), .OUT(n5479) );
  NAND2 U4026 ( .A(n5479), .B(n1766), .OUT(n4429) );
  NAND2 U4027 ( .A(n3292), .B(n4429), .OUT(n1877) );
  NAND2 U4028 ( .A(\mult_49/ab[26][3] ), .B(n1767), .OUT(n1876) );
  INV U4029 ( .IN(n1875), .OUT(n5480) );
  NAND2 U4030 ( .A(n5480), .B(n1874), .OUT(n4506) );
  NAND2 U4031 ( .A(n3373), .B(n4506), .OUT(n4803) );
  NAND2 U4032 ( .A(\mult_49/ab[27][3] ), .B(n1875), .OUT(n4507) );
  NAND2 U4033 ( .A(n5133), .B(n431), .OUT(n3799) );
  NAND2 U4034 ( .A(n2264), .B(n3799), .OUT(n513) );
  NAND2 U4035 ( .A(\mult_49/ab[9][2] ), .B(n432), .OUT(n512) );
  INV U4036 ( .IN(n511), .OUT(n5481) );
  NAND2 U4037 ( .A(n5481), .B(n546), .OUT(n4509) );
  NAND2 U4038 ( .A(n2377), .B(n4509), .OUT(n549) );
  NAND2 U4039 ( .A(\mult_49/ab[10][2] ), .B(n511), .OUT(n548) );
  INV U4040 ( .IN(n547), .OUT(n5482) );
  NAND2 U4041 ( .A(n5482), .B(n586), .OUT(n4511) );
  NAND2 U4042 ( .A(n2407), .B(n4511), .OUT(n589) );
  NAND2 U4043 ( .A(\mult_49/ab[11][2] ), .B(n547), .OUT(n588) );
  INV U4044 ( .IN(n587), .OUT(n5483) );
  NAND2 U4045 ( .A(n5483), .B(n630), .OUT(n4513) );
  NAND2 U4046 ( .A(n2440), .B(n4513), .OUT(n633) );
  NAND2 U4047 ( .A(\mult_49/ab[12][2] ), .B(n587), .OUT(n632) );
  INV U4048 ( .IN(n631), .OUT(n5484) );
  NAND2 U4049 ( .A(n5484), .B(n678), .OUT(n4515) );
  NAND2 U4050 ( .A(n2476), .B(n4515), .OUT(n681) );
  NAND2 U4051 ( .A(\mult_49/ab[13][2] ), .B(n631), .OUT(n680) );
  INV U4052 ( .IN(n679), .OUT(n5485) );
  NAND2 U4053 ( .A(n5485), .B(n730), .OUT(n4517) );
  NAND2 U4054 ( .A(n2515), .B(n4517), .OUT(n733) );
  NAND2 U4055 ( .A(\mult_49/ab[14][2] ), .B(n679), .OUT(n732) );
  INV U4056 ( .IN(n731), .OUT(n5486) );
  NAND2 U4057 ( .A(n5486), .B(n786), .OUT(n4519) );
  NAND2 U4058 ( .A(n2557), .B(n4519), .OUT(n789) );
  NAND2 U4059 ( .A(\mult_49/ab[15][2] ), .B(n731), .OUT(n788) );
  INV U4060 ( .IN(n787), .OUT(n5487) );
  NAND2 U4061 ( .A(n5487), .B(n846), .OUT(n4521) );
  NAND2 U4062 ( .A(n2602), .B(n4521), .OUT(n849) );
  NAND2 U4063 ( .A(\mult_49/ab[16][2] ), .B(n787), .OUT(n848) );
  INV U4064 ( .IN(n847), .OUT(n5488) );
  NAND2 U4065 ( .A(n5488), .B(n910), .OUT(n4523) );
  NAND2 U4066 ( .A(n2650), .B(n4523), .OUT(n913) );
  NAND2 U4067 ( .A(\mult_49/ab[17][2] ), .B(n847), .OUT(n912) );
  INV U4068 ( .IN(n911), .OUT(n5489) );
  NAND2 U4069 ( .A(n5489), .B(n978), .OUT(n4525) );
  NAND2 U4070 ( .A(n2701), .B(n4525), .OUT(n981) );
  NAND2 U4071 ( .A(\mult_49/ab[18][2] ), .B(n911), .OUT(n980) );
  INV U4072 ( .IN(n979), .OUT(n5490) );
  NAND2 U4073 ( .A(n5490), .B(n1050), .OUT(n4527) );
  NAND2 U4074 ( .A(n2755), .B(n4527), .OUT(n1053) );
  NAND2 U4075 ( .A(\mult_49/ab[19][2] ), .B(n979), .OUT(n1052) );
  INV U4076 ( .IN(n1051), .OUT(n5491) );
  NAND2 U4077 ( .A(n5491), .B(n1126), .OUT(n4529) );
  NAND2 U4078 ( .A(n2812), .B(n4529), .OUT(n1129) );
  NAND2 U4079 ( .A(\mult_49/ab[20][2] ), .B(n1051), .OUT(n1128) );
  INV U4080 ( .IN(n1127), .OUT(n5492) );
  NAND2 U4081 ( .A(n5492), .B(n1206), .OUT(n4531) );
  NAND2 U4082 ( .A(n2872), .B(n4531), .OUT(n1209) );
  NAND2 U4083 ( .A(\mult_49/ab[21][2] ), .B(n1127), .OUT(n1208) );
  INV U4084 ( .IN(n1207), .OUT(n5493) );
  NAND2 U4085 ( .A(n5493), .B(n1290), .OUT(n4533) );
  NAND2 U4086 ( .A(n2935), .B(n4533), .OUT(n1293) );
  NAND2 U4087 ( .A(\mult_49/ab[22][2] ), .B(n1207), .OUT(n1292) );
  INV U4088 ( .IN(n1291), .OUT(n5494) );
  NAND2 U4089 ( .A(n5494), .B(n1378), .OUT(n4535) );
  NAND2 U4090 ( .A(n3001), .B(n4535), .OUT(n1381) );
  NAND2 U4091 ( .A(\mult_49/ab[23][2] ), .B(n1291), .OUT(n1380) );
  INV U4092 ( .IN(n1379), .OUT(n5495) );
  NAND2 U4093 ( .A(n5495), .B(n1470), .OUT(n4537) );
  NAND2 U4094 ( .A(n3070), .B(n4537), .OUT(n1473) );
  NAND2 U4095 ( .A(\mult_49/ab[24][2] ), .B(n1379), .OUT(n1472) );
  INV U4096 ( .IN(n1471), .OUT(n5496) );
  NAND2 U4097 ( .A(n5496), .B(n1566), .OUT(n4539) );
  NAND2 U4098 ( .A(n3142), .B(n4539), .OUT(n1569) );
  NAND2 U4099 ( .A(\mult_49/ab[25][2] ), .B(n1471), .OUT(n1568) );
  INV U4100 ( .IN(n1567), .OUT(n5497) );
  NAND2 U4101 ( .A(n5497), .B(n1666), .OUT(n4541) );
  NAND2 U4102 ( .A(n3217), .B(n4541), .OUT(n1669) );
  NAND2 U4103 ( .A(\mult_49/ab[26][2] ), .B(n1567), .OUT(n1668) );
  INV U4104 ( .IN(n1667), .OUT(n5498) );
  NAND2 U4105 ( .A(n5498), .B(n1770), .OUT(n4543) );
  NAND2 U4106 ( .A(n3295), .B(n4543), .OUT(n1773) );
  NAND2 U4107 ( .A(\mult_49/ab[27][2] ), .B(n1667), .OUT(n1772) );
  INV U4108 ( .IN(n1771), .OUT(n5499) );
  NAND2 U4109 ( .A(n5499), .B(n1878), .OUT(n4545) );
  NAND2 U4110 ( .A(n3376), .B(n4545), .OUT(n4851) );
  NAND2 U4111 ( .A(\mult_49/ab[28][2] ), .B(n1771), .OUT(n4546) );
  NAND2 U4112 ( .A(n5142), .B(n467), .OUT(n3801) );
  NAND2 U4113 ( .A(n2288), .B(n3801), .OUT(n1881) );
  NAND2 U4114 ( .A(\mult_49/ab[10][1] ), .B(n468), .OUT(n1880) );
  INV U4115 ( .IN(n1879), .OUT(n5500) );
  NAND2 U4116 ( .A(n5500), .B(n1882), .OUT(n4548) );
  NAND2 U4117 ( .A(n3406), .B(n4548), .OUT(n1885) );
  NAND2 U4118 ( .A(\mult_49/ab[11][1] ), .B(n1879), .OUT(n1884) );
  INV U4119 ( .IN(n1883), .OUT(n5501) );
  NAND2 U4120 ( .A(n5501), .B(n1886), .OUT(n4550) );
  NAND2 U4121 ( .A(n3412), .B(n4550), .OUT(n1889) );
  NAND2 U4122 ( .A(\mult_49/ab[12][1] ), .B(n1883), .OUT(n1888) );
  INV U4123 ( .IN(n1887), .OUT(n5502) );
  NAND2 U4124 ( .A(n5502), .B(n1890), .OUT(n4552) );
  NAND2 U4125 ( .A(n3418), .B(n4552), .OUT(n1893) );
  NAND2 U4126 ( .A(\mult_49/ab[13][1] ), .B(n1887), .OUT(n1892) );
  INV U4127 ( .IN(n1891), .OUT(n5503) );
  NAND2 U4128 ( .A(n5503), .B(n1894), .OUT(n4554) );
  NAND2 U4129 ( .A(n3424), .B(n4554), .OUT(n1897) );
  NAND2 U4130 ( .A(\mult_49/ab[14][1] ), .B(n1891), .OUT(n1896) );
  INV U4131 ( .IN(n1895), .OUT(n5504) );
  NAND2 U4132 ( .A(n5504), .B(n1898), .OUT(n4556) );
  NAND2 U4133 ( .A(n3430), .B(n4556), .OUT(n1901) );
  NAND2 U4134 ( .A(\mult_49/ab[15][1] ), .B(n1895), .OUT(n1900) );
  INV U4135 ( .IN(n1899), .OUT(n5505) );
  NAND2 U4136 ( .A(n5505), .B(n1902), .OUT(n4558) );
  NAND2 U4137 ( .A(n3436), .B(n4558), .OUT(n1905) );
  NAND2 U4138 ( .A(\mult_49/ab[16][1] ), .B(n1899), .OUT(n1904) );
  INV U4139 ( .IN(n1903), .OUT(n5506) );
  NAND2 U4140 ( .A(n5506), .B(n1906), .OUT(n4560) );
  NAND2 U4141 ( .A(n3442), .B(n4560), .OUT(n1909) );
  NAND2 U4142 ( .A(\mult_49/ab[17][1] ), .B(n1903), .OUT(n1908) );
  INV U4143 ( .IN(n1907), .OUT(n5507) );
  NAND2 U4144 ( .A(n5507), .B(n1910), .OUT(n4562) );
  NAND2 U4145 ( .A(n3448), .B(n4562), .OUT(n1913) );
  NAND2 U4146 ( .A(\mult_49/ab[18][1] ), .B(n1907), .OUT(n1912) );
  INV U4147 ( .IN(n1911), .OUT(n5508) );
  NAND2 U4148 ( .A(n5508), .B(n1914), .OUT(n4564) );
  NAND2 U4149 ( .A(n3454), .B(n4564), .OUT(n1917) );
  NAND2 U4150 ( .A(\mult_49/ab[19][1] ), .B(n1911), .OUT(n1916) );
  INV U4151 ( .IN(n1915), .OUT(n5509) );
  NAND2 U4152 ( .A(n5509), .B(n1918), .OUT(n4566) );
  NAND2 U4153 ( .A(n3460), .B(n4566), .OUT(n1921) );
  NAND2 U4154 ( .A(\mult_49/ab[20][1] ), .B(n1915), .OUT(n1920) );
  INV U4155 ( .IN(n1919), .OUT(n5510) );
  NAND2 U4156 ( .A(n5510), .B(n1922), .OUT(n4568) );
  NAND2 U4157 ( .A(n3466), .B(n4568), .OUT(n1925) );
  NAND2 U4158 ( .A(\mult_49/ab[21][1] ), .B(n1919), .OUT(n1924) );
  INV U4159 ( .IN(n1923), .OUT(n5511) );
  NAND2 U4160 ( .A(n5511), .B(n1926), .OUT(n4570) );
  NAND2 U4161 ( .A(n3472), .B(n4570), .OUT(n1929) );
  NAND2 U4162 ( .A(\mult_49/ab[22][1] ), .B(n1923), .OUT(n1928) );
  INV U4163 ( .IN(n1927), .OUT(n5512) );
  NAND2 U4164 ( .A(n5512), .B(n1930), .OUT(n4572) );
  NAND2 U4165 ( .A(n3478), .B(n4572), .OUT(n1933) );
  NAND2 U4166 ( .A(\mult_49/ab[23][1] ), .B(n1927), .OUT(n1932) );
  INV U4167 ( .IN(n1931), .OUT(n5513) );
  NAND2 U4168 ( .A(n5513), .B(n1934), .OUT(n4574) );
  NAND2 U4169 ( .A(n3484), .B(n4574), .OUT(n1937) );
  NAND2 U4170 ( .A(\mult_49/ab[24][1] ), .B(n1931), .OUT(n1936) );
  INV U4171 ( .IN(n1935), .OUT(n5514) );
  NAND2 U4172 ( .A(n5514), .B(n1938), .OUT(n4576) );
  NAND2 U4173 ( .A(n3490), .B(n4576), .OUT(n1941) );
  NAND2 U4174 ( .A(\mult_49/ab[25][1] ), .B(n1935), .OUT(n1940) );
  INV U4175 ( .IN(n1939), .OUT(n5515) );
  NAND2 U4176 ( .A(n5515), .B(n1942), .OUT(n4578) );
  NAND2 U4177 ( .A(n3496), .B(n4578), .OUT(n1945) );
  NAND2 U4178 ( .A(\mult_49/ab[26][1] ), .B(n1939), .OUT(n1944) );
  INV U4179 ( .IN(n1943), .OUT(n5516) );
  NAND2 U4180 ( .A(n5516), .B(n1946), .OUT(n4580) );
  NAND2 U4181 ( .A(n3502), .B(n4580), .OUT(n1949) );
  NAND2 U4182 ( .A(\mult_49/ab[27][1] ), .B(n1943), .OUT(n1948) );
  INV U4183 ( .IN(n1947), .OUT(n5517) );
  NAND2 U4184 ( .A(n5517), .B(n1950), .OUT(n4582) );
  NAND2 U4185 ( .A(n3508), .B(n4582), .OUT(n1953) );
  NAND2 U4186 ( .A(\mult_49/ab[28][1] ), .B(n1947), .OUT(n1952) );
  INV U4187 ( .IN(n1951), .OUT(n5518) );
  NAND2 U4188 ( .A(n5518), .B(n1954), .OUT(n4584) );
  NAND2 U4189 ( .A(n3514), .B(n4584), .OUT(n4847) );
  NAND2 U4190 ( .A(\mult_49/ab[29][1] ), .B(n1951), .OUT(n4585) );
  NAND2 U4191 ( .A(n5155), .B(n507), .OUT(n3803) );
  NAND2 U4192 ( .A(n5519), .B(n3803), .OUT(n1957) );
  NAND2 U4193 ( .A(\mult_49/ab[11][0] ), .B(n508), .OUT(n1956) );
  INV U4194 ( .IN(n1955), .OUT(n5520) );
  NAND2 U4195 ( .A(n3409), .B(n4776), .OUT(n1961) );
  INV U4196 ( .IN(n1959), .OUT(n5521) );
  NAND2 U4197 ( .A(n5522), .B(n4774), .OUT(n1965) );
  INV U4198 ( .IN(n1963), .OUT(n5523) );
  NAND2 U4199 ( .A(n3421), .B(n4772), .OUT(n1969) );
  INV U4200 ( .IN(n1967), .OUT(n5524) );
  NAND2 U4201 ( .A(n5525), .B(n4770), .OUT(n1973) );
  INV U4202 ( .IN(n1971), .OUT(n5526) );
  NAND2 U4203 ( .A(n3433), .B(n4768), .OUT(n1977) );
  INV U4204 ( .IN(n1975), .OUT(n5527) );
  NAND2 U4205 ( .A(n5528), .B(n4766), .OUT(n1981) );
  INV U4206 ( .IN(n1979), .OUT(n5529) );
  NAND2 U4207 ( .A(n3445), .B(n4764), .OUT(n1985) );
  INV U4208 ( .IN(n1983), .OUT(n5530) );
  NAND2 U4209 ( .A(n5531), .B(n4762), .OUT(n1989) );
  INV U4210 ( .IN(n1987), .OUT(n5532) );
  NAND2 U4211 ( .A(n3457), .B(n4760), .OUT(n1993) );
  INV U4212 ( .IN(n1991), .OUT(n5533) );
  NAND2 U4213 ( .A(n5534), .B(n4758), .OUT(n1997) );
  INV U4214 ( .IN(n1995), .OUT(n5535) );
  NAND2 U4215 ( .A(n3469), .B(n4754), .OUT(n2001) );
  INV U4216 ( .IN(n1999), .OUT(n5536) );
  NAND2 U4217 ( .A(n5537), .B(n4752), .OUT(n2005) );
  INV U4218 ( .IN(n2003), .OUT(n5538) );
  NAND2 U4219 ( .A(n3481), .B(n4750), .OUT(n2009) );
  INV U4220 ( .IN(n2007), .OUT(n5539) );
  NAND2 U4221 ( .A(n5540), .B(n4748), .OUT(n2013) );
  INV U4222 ( .IN(n2011), .OUT(n5541) );
  NAND2 U4223 ( .A(n3493), .B(n4746), .OUT(n2017) );
  INV U4224 ( .IN(n2015), .OUT(n5542) );
  NAND2 U4225 ( .A(n5543), .B(n4744), .OUT(n2021) );
  INV U4226 ( .IN(n2019), .OUT(n5544) );
  NAND2 U4227 ( .A(n3505), .B(n4742), .OUT(n2025) );
  INV U4228 ( .IN(n2023), .OUT(n5545) );
  NAND2 U4229 ( .A(n5546), .B(n4740), .OUT(n2029) );
  INV U4230 ( .IN(n2027), .OUT(n5547) );
  NAND2 U4231 ( .A(n3517), .B(n4737), .OUT(n4849) );
  NAND2 U4232 ( .A(n2069), .B(n2070), .OUT(n5548) );
  NAND2 U4233 ( .A(n2091), .B(n5548), .OUT(n4912) );
  NAND2 U4234 ( .A(B[1]), .B(A[1]), .OUT(n4911) );
  NAND2 U4235 ( .A(n2047), .B(n2048), .OUT(n5549) );
  NAND2 U4236 ( .A(n5549), .B(n4910), .OUT(n4906) );
  NAND2 U4237 ( .A(B[2]), .B(A[2]), .OUT(n4905) );
  NAND2 U4238 ( .A(n2043), .B(n2044), .OUT(n5550) );
  NAND2 U4239 ( .A(n5550), .B(n4904), .OUT(n4900) );
  NAND2 U4240 ( .A(B[3]), .B(A[3]), .OUT(n4899) );
  NAND2 U4241 ( .A(n2041), .B(n2042), .OUT(n5551) );
  NAND2 U4242 ( .A(n5551), .B(n4898), .OUT(n4894) );
  NAND2 U4243 ( .A(B[4]), .B(A[4]), .OUT(n4893) );
  NAND2 U4244 ( .A(n2039), .B(n2040), .OUT(n5552) );
  NAND2 U4245 ( .A(n5552), .B(n4892), .OUT(n4888) );
  NAND2 U4246 ( .A(B[5]), .B(A[5]), .OUT(n4887) );
  INV U4247 ( .IN(n2092), .OUT(n289) );
  NAND2 U4248 ( .A(A[0]), .B(\mult_49/B_notx[0] ), .OUT(n290) );
  NAND2 U4249 ( .A(n2092), .B(B[1]), .OUT(n5553) );
  NAND2 U4250 ( .A(A[1]), .B(n5553), .OUT(n2095) );
  NAND2 U4251 ( .A(n289), .B(n2070), .OUT(n2094) );
  INV U4252 ( .IN(n2093), .OUT(n5554) );
  NAND2 U4253 ( .A(n5554), .B(B[2]), .OUT(n5555) );
  NAND2 U4254 ( .A(A[2]), .B(n5555), .OUT(n2098) );
  NAND2 U4255 ( .A(n2093), .B(n2048), .OUT(n2097) );
  INV U4256 ( .IN(n2096), .OUT(n5556) );
  NAND2 U4257 ( .A(n5556), .B(B[3]), .OUT(n5557) );
  NAND2 U4258 ( .A(A[3]), .B(n5557), .OUT(n2101) );
  NAND2 U4259 ( .A(n2096), .B(n2044), .OUT(n2100) );
  INV U4260 ( .IN(n2099), .OUT(n5558) );
  NAND2 U4261 ( .A(n5558), .B(B[4]), .OUT(n5559) );
  NAND2 U4262 ( .A(A[4]), .B(n5559), .OUT(n2104) );
  NAND2 U4263 ( .A(n2099), .B(n2042), .OUT(n2103) );
  INV U4264 ( .IN(n2102), .OUT(n5560) );
  NAND2 U4265 ( .A(n5560), .B(B[5]), .OUT(n5561) );
  NAND2 U4266 ( .A(A[5]), .B(n5561), .OUT(n2107) );
  NAND2 U4267 ( .A(n2102), .B(n2040), .OUT(n2106) );
  INV U4268 ( .IN(n2105), .OUT(n5562) );
  NAND2 U4269 ( .A(n5562), .B(B[6]), .OUT(n5563) );
  NAND2 U4270 ( .A(A[6]), .B(n5563), .OUT(n2110) );
  NAND2 U4271 ( .A(n2105), .B(n2038), .OUT(n2109) );
  INV U4272 ( .IN(n2108), .OUT(n5564) );
  NAND2 U4273 ( .A(n5564), .B(B[7]), .OUT(n5565) );
  NAND2 U4274 ( .A(A[7]), .B(n5565), .OUT(n2113) );
  NAND2 U4275 ( .A(n2108), .B(n2036), .OUT(n2112) );
  INV U4276 ( .IN(n2111), .OUT(n5566) );
  NAND2 U4277 ( .A(n5566), .B(B[8]), .OUT(n5567) );
  NAND2 U4278 ( .A(A[8]), .B(n5567), .OUT(n2116) );
  NAND2 U4279 ( .A(n2111), .B(n2034), .OUT(n2115) );
  INV U4280 ( .IN(n2114), .OUT(n5568) );
  NAND2 U4281 ( .A(n5568), .B(B[9]), .OUT(n5569) );
  NAND2 U4282 ( .A(A[9]), .B(n5569), .OUT(n2119) );
  NAND2 U4283 ( .A(n2114), .B(n2032), .OUT(n2118) );
  INV U4284 ( .IN(n2117), .OUT(n5570) );
  NAND2 U4285 ( .A(n5570), .B(B[10]), .OUT(n5571) );
  NAND2 U4286 ( .A(A[10]), .B(n5571), .OUT(n2122) );
  NAND2 U4287 ( .A(n2117), .B(n2090), .OUT(n2121) );
  INV U4288 ( .IN(n2120), .OUT(n5572) );
  NAND2 U4289 ( .A(n5572), .B(B[11]), .OUT(n5573) );
  NAND2 U4290 ( .A(A[11]), .B(n5573), .OUT(n2125) );
  NAND2 U4291 ( .A(n2120), .B(n2088), .OUT(n2124) );
  INV U4292 ( .IN(n2123), .OUT(n5574) );
  NAND2 U4293 ( .A(n5574), .B(B[12]), .OUT(n5575) );
  NAND2 U4294 ( .A(A[12]), .B(n5575), .OUT(n2128) );
  NAND2 U4295 ( .A(n2123), .B(n2086), .OUT(n2127) );
  INV U4296 ( .IN(n2126), .OUT(n5576) );
  NAND2 U4297 ( .A(n5576), .B(B[13]), .OUT(n5577) );
  NAND2 U4298 ( .A(A[13]), .B(n5577), .OUT(n2131) );
  NAND2 U4299 ( .A(n2126), .B(n2084), .OUT(n2130) );
  INV U4300 ( .IN(n2129), .OUT(n5578) );
  NAND2 U4301 ( .A(n5578), .B(B[14]), .OUT(n5579) );
  NAND2 U4302 ( .A(A[14]), .B(n5579), .OUT(n2134) );
  NAND2 U4303 ( .A(n2129), .B(n2082), .OUT(n2133) );
  INV U4304 ( .IN(n2132), .OUT(n5580) );
  NAND2 U4305 ( .A(n5580), .B(B[15]), .OUT(n5581) );
  NAND2 U4306 ( .A(A[15]), .B(n5581), .OUT(n2137) );
  NAND2 U4307 ( .A(n2132), .B(n2080), .OUT(n2136) );
  INV U4308 ( .IN(n2135), .OUT(n5582) );
  NAND2 U4309 ( .A(n5582), .B(B[16]), .OUT(n5583) );
  NAND2 U4310 ( .A(A[16]), .B(n5583), .OUT(n2140) );
  NAND2 U4311 ( .A(n2135), .B(n2078), .OUT(n2139) );
  INV U4312 ( .IN(n2138), .OUT(n5584) );
  NAND2 U4313 ( .A(n5584), .B(B[17]), .OUT(n5585) );
  NAND2 U4314 ( .A(A[17]), .B(n5585), .OUT(n2143) );
  NAND2 U4315 ( .A(n2138), .B(n2076), .OUT(n2142) );
  INV U4316 ( .IN(n2141), .OUT(n5586) );
  NAND2 U4317 ( .A(n5586), .B(B[18]), .OUT(n5587) );
  NAND2 U4318 ( .A(A[18]), .B(n5587), .OUT(n2146) );
  NAND2 U4319 ( .A(n2141), .B(n2074), .OUT(n2145) );
  INV U4320 ( .IN(n2144), .OUT(n5588) );
  NAND2 U4321 ( .A(n5588), .B(B[19]), .OUT(n5589) );
  NAND2 U4322 ( .A(A[19]), .B(n5589), .OUT(n2149) );
  NAND2 U4323 ( .A(n2144), .B(n2072), .OUT(n2148) );
  INV U4324 ( .IN(n2147), .OUT(n5590) );
  NAND2 U4325 ( .A(n5590), .B(B[20]), .OUT(n5591) );
  NAND2 U4326 ( .A(A[20]), .B(n5591), .OUT(n2152) );
  NAND2 U4327 ( .A(n2147), .B(n2068), .OUT(n2151) );
  INV U4328 ( .IN(n2150), .OUT(n5592) );
  NAND2 U4329 ( .A(n5592), .B(B[21]), .OUT(n5593) );
  NAND2 U4330 ( .A(A[21]), .B(n5593), .OUT(n2155) );
  NAND2 U4331 ( .A(n2150), .B(n2066), .OUT(n2154) );
  INV U4332 ( .IN(n2153), .OUT(n5594) );
  NAND2 U4333 ( .A(n5594), .B(B[22]), .OUT(n5595) );
  NAND2 U4334 ( .A(A[22]), .B(n5595), .OUT(n2158) );
  NAND2 U4335 ( .A(n2153), .B(n2064), .OUT(n2157) );
  INV U4336 ( .IN(n2156), .OUT(n5596) );
  NAND2 U4337 ( .A(n5596), .B(B[23]), .OUT(n5597) );
  NAND2 U4338 ( .A(A[23]), .B(n5597), .OUT(n2161) );
  NAND2 U4339 ( .A(n2156), .B(n2062), .OUT(n2160) );
  INV U4340 ( .IN(n2159), .OUT(n5598) );
  NAND2 U4341 ( .A(n5598), .B(B[24]), .OUT(n5599) );
  NAND2 U4342 ( .A(A[24]), .B(n5599), .OUT(n2164) );
  NAND2 U4343 ( .A(n2159), .B(n2060), .OUT(n2163) );
  INV U4344 ( .IN(n2162), .OUT(n5600) );
  NAND2 U4345 ( .A(n5600), .B(B[25]), .OUT(n5601) );
  NAND2 U4346 ( .A(A[25]), .B(n5601), .OUT(n2167) );
  NAND2 U4347 ( .A(n2162), .B(n2058), .OUT(n2166) );
  INV U4348 ( .IN(n2165), .OUT(n5602) );
  NAND2 U4349 ( .A(n5602), .B(B[26]), .OUT(n5603) );
  NAND2 U4350 ( .A(A[26]), .B(n5603), .OUT(n2170) );
  NAND2 U4351 ( .A(n2165), .B(n2056), .OUT(n2169) );
  INV U4352 ( .IN(n2168), .OUT(n5604) );
  NAND2 U4353 ( .A(n5604), .B(B[27]), .OUT(n5605) );
  NAND2 U4354 ( .A(A[27]), .B(n5605), .OUT(n2173) );
  NAND2 U4355 ( .A(n2168), .B(n2054), .OUT(n2172) );
  INV U4356 ( .IN(n2171), .OUT(n5606) );
  NAND2 U4357 ( .A(n5606), .B(B[28]), .OUT(n5607) );
  NAND2 U4358 ( .A(A[28]), .B(n5607), .OUT(n2176) );
  NAND2 U4359 ( .A(n2171), .B(n2052), .OUT(n2175) );
  INV U4360 ( .IN(n2174), .OUT(n5608) );
  NAND2 U4361 ( .A(n5608), .B(B[29]), .OUT(n5609) );
  NAND2 U4362 ( .A(A[29]), .B(n5609), .OUT(n2179) );
  NAND2 U4363 ( .A(n2174), .B(n2050), .OUT(n2178) );
  INV U4364 ( .IN(n2177), .OUT(n5610) );
  NAND2 U4365 ( .A(n5610), .B(B[30]), .OUT(n5611) );
  NAND2 U4366 ( .A(A[30]), .B(n5611), .OUT(n4918) );
  NAND2 U4367 ( .A(n2177), .B(n2046), .OUT(n4917) );
  NAND2 U4368 ( .A(n2037), .B(n2038), .OUT(n5612) );
  NAND2 U4369 ( .A(n5612), .B(n4886), .OUT(n5066) );
  NAND2 U4370 ( .A(B[6]), .B(A[6]), .OUT(n5065) );
  NAND2 U4371 ( .A(n2035), .B(n2036), .OUT(n5613) );
  NAND2 U4372 ( .A(n5613), .B(n5064), .OUT(n5060) );
  NAND2 U4373 ( .A(B[7]), .B(A[7]), .OUT(n5059) );
  NAND2 U4374 ( .A(n2033), .B(n2034), .OUT(n5614) );
  NAND2 U4375 ( .A(n5614), .B(n5058), .OUT(n5054) );
  NAND2 U4376 ( .A(B[8]), .B(A[8]), .OUT(n5053) );
  NAND2 U4377 ( .A(n2031), .B(n2032), .OUT(n5615) );
  NAND2 U4378 ( .A(n5615), .B(n5052), .OUT(n5048) );
  NAND2 U4379 ( .A(B[9]), .B(A[9]), .OUT(n5047) );
  NAND2 U4380 ( .A(n2089), .B(n2090), .OUT(n5616) );
  NAND2 U4381 ( .A(n5616), .B(n5046), .OUT(n5042) );
  NAND2 U4382 ( .A(B[10]), .B(A[10]), .OUT(n5041) );
  NAND2 U4383 ( .A(n2087), .B(n2088), .OUT(n5617) );
  NAND2 U4384 ( .A(n5617), .B(n5040), .OUT(n5036) );
  NAND2 U4385 ( .A(B[11]), .B(A[11]), .OUT(n5035) );
  NAND2 U4386 ( .A(n2085), .B(n2086), .OUT(n5618) );
  NAND2 U4387 ( .A(n5618), .B(n5034), .OUT(n5030) );
  NAND2 U4388 ( .A(B[12]), .B(A[12]), .OUT(n5029) );
  NAND2 U4389 ( .A(n2083), .B(n2084), .OUT(n5619) );
  NAND2 U4390 ( .A(n5619), .B(n5028), .OUT(n5024) );
  NAND2 U4391 ( .A(B[13]), .B(A[13]), .OUT(n5023) );
  NAND2 U4392 ( .A(n2081), .B(n2082), .OUT(n5620) );
  NAND2 U4393 ( .A(n5620), .B(n5022), .OUT(n5018) );
  NAND2 U4394 ( .A(B[14]), .B(A[14]), .OUT(n5017) );
  NAND2 U4395 ( .A(n2079), .B(n2080), .OUT(n5621) );
  NAND2 U4396 ( .A(n5621), .B(n5016), .OUT(n5012) );
  NAND2 U4397 ( .A(B[15]), .B(A[15]), .OUT(n5011) );
  NAND2 U4398 ( .A(n2077), .B(n2078), .OUT(n5622) );
  NAND2 U4399 ( .A(n5622), .B(n5010), .OUT(n5006) );
  NAND2 U4400 ( .A(B[16]), .B(A[16]), .OUT(n5005) );
  NAND2 U4401 ( .A(n2075), .B(n2076), .OUT(n5623) );
  NAND2 U4402 ( .A(n5623), .B(n5004), .OUT(n5000) );
  NAND2 U4403 ( .A(B[17]), .B(A[17]), .OUT(n4999) );
  NAND2 U4404 ( .A(n2073), .B(n2074), .OUT(n5624) );
  NAND2 U4405 ( .A(n5624), .B(n4998), .OUT(n4994) );
  NAND2 U4406 ( .A(B[18]), .B(A[18]), .OUT(n4993) );
  NAND2 U4407 ( .A(n2071), .B(n2072), .OUT(n5625) );
  NAND2 U4408 ( .A(n5625), .B(n4992), .OUT(n4988) );
  NAND2 U4409 ( .A(B[19]), .B(A[19]), .OUT(n4987) );
  NAND2 U4410 ( .A(n2067), .B(n2068), .OUT(n5626) );
  NAND2 U4411 ( .A(n5626), .B(n4986), .OUT(n4982) );
  NAND2 U4412 ( .A(B[20]), .B(A[20]), .OUT(n4981) );
  NAND2 U4413 ( .A(n2065), .B(n2066), .OUT(n5627) );
  NAND2 U4414 ( .A(n5627), .B(n4980), .OUT(n4976) );
  NAND2 U4415 ( .A(B[21]), .B(A[21]), .OUT(n4975) );
  NAND2 U4416 ( .A(n2063), .B(n2064), .OUT(n5628) );
  NAND2 U4417 ( .A(n5628), .B(n4974), .OUT(n4970) );
  NAND2 U4418 ( .A(B[22]), .B(A[22]), .OUT(n4969) );
  NAND2 U4419 ( .A(n2061), .B(n2062), .OUT(n5629) );
  NAND2 U4420 ( .A(n5629), .B(n4968), .OUT(n4964) );
  NAND2 U4421 ( .A(B[23]), .B(A[23]), .OUT(n4963) );
  NAND2 U4422 ( .A(n2059), .B(n2060), .OUT(n5630) );
  NAND2 U4423 ( .A(n5630), .B(n4962), .OUT(n4958) );
  NAND2 U4424 ( .A(B[24]), .B(A[24]), .OUT(n4957) );
  NAND2 U4425 ( .A(n2057), .B(n2058), .OUT(n5631) );
  NAND2 U4426 ( .A(n5631), .B(n4956), .OUT(n4952) );
  NAND2 U4427 ( .A(B[25]), .B(A[25]), .OUT(n4951) );
  NAND2 U4428 ( .A(n2055), .B(n2056), .OUT(n5632) );
  NAND2 U4429 ( .A(n5632), .B(n4950), .OUT(n4946) );
  NAND2 U4430 ( .A(B[26]), .B(A[26]), .OUT(n4945) );
  NAND2 U4431 ( .A(n2053), .B(n2054), .OUT(n5633) );
  NAND2 U4432 ( .A(n5633), .B(n4944), .OUT(n4940) );
  NAND2 U4433 ( .A(B[27]), .B(A[27]), .OUT(n4939) );
  NAND2 U4434 ( .A(n2051), .B(n2052), .OUT(n5634) );
  NAND2 U4435 ( .A(n5634), .B(n4938), .OUT(n4934) );
  NAND2 U4436 ( .A(B[28]), .B(A[28]), .OUT(n4933) );
  NAND2 U4437 ( .A(n2049), .B(n2050), .OUT(n5635) );
  NAND2 U4438 ( .A(n5635), .B(n4932), .OUT(n4928) );
  NAND2 U4439 ( .A(B[29]), .B(A[29]), .OUT(n4927) );
  NAND2 U4440 ( .A(n2045), .B(n2046), .OUT(n5636) );
  NAND2 U4441 ( .A(n5636), .B(n4926), .OUT(n4921) );
  NAND2 U4442 ( .A(B[30]), .B(A[30]), .OUT(n4920) );
  NAND2 U4443 ( .A(\mult_49/ab[0][11] ), .B(n515), .OUT(n2182) );
  NAND2 U4444 ( .A(\mult_49/ab[1][10] ), .B(n516), .OUT(n2181) );
  NAND2 U4445 ( .A(n291), .B(n294), .OUT(n3785) );
  NAND2 U4446 ( .A(\mult_49/ab[2][9] ), .B(n5089), .OUT(n3784) );
  NAND2 U4447 ( .A(n2180), .B(n5637), .OUT(n2185) );
  NOR2 U4448 ( .A(n5637), .B(n2180), .OUT(n5638) );
  NAND2 U4449 ( .A(\mult_49/ab[0][10] ), .B(n293), .OUT(n2188) );
  NAND2 U4450 ( .A(\mult_49/ab[1][9] ), .B(n292), .OUT(n2187) );
  NOR2 U4451 ( .A(n5639), .B(n3786), .OUT(n2191) );
  NOR2 U4452 ( .A(n5640), .B(n2183), .OUT(n2190) );
  NAND2 U4453 ( .A(\mult_49/ab[0][9] ), .B(n298), .OUT(n2194) );
  NAND2 U4454 ( .A(\mult_49/ab[1][8] ), .B(n297), .OUT(n2193) );
  NAND2 U4455 ( .A(n296), .B(n295), .OUT(n3768) );
  NAND2 U4456 ( .A(\mult_49/ab[2][8] ), .B(n5090), .OUT(n3767) );
  NAND2 U4457 ( .A(n2186), .B(n5641), .OUT(n2197) );
  NOR2 U4458 ( .A(n5641), .B(n2186), .OUT(n5642) );
  NOR2 U4459 ( .A(n2189), .B(n3788), .OUT(n5643) );
  NAND2 U4460 ( .A(n3788), .B(n2189), .OUT(n2199) );
  NAND2 U4461 ( .A(\mult_49/ab[0][8] ), .B(n306), .OUT(n2203) );
  NAND2 U4462 ( .A(\mult_49/ab[1][7] ), .B(n305), .OUT(n2202) );
  NAND2 U4463 ( .A(n304), .B(n303), .OUT(n3753) );
  NAND2 U4464 ( .A(\mult_49/ab[2][7] ), .B(n5091), .OUT(n3752) );
  NAND2 U4465 ( .A(n2192), .B(n5644), .OUT(n2206) );
  NOR2 U4466 ( .A(n5644), .B(n2192), .OUT(n5645) );
  NOR2 U4467 ( .A(n5646), .B(n3769), .OUT(n2209) );
  NOR2 U4468 ( .A(n5647), .B(n2195), .OUT(n2208) );
  NAND2 U4469 ( .A(n2198), .B(n5649), .OUT(n5648) );
  NOR2 U4470 ( .A(n5649), .B(n2198), .OUT(n2211) );
  NAND2 U4471 ( .A(\mult_49/ab[0][7] ), .B(n318), .OUT(n2215) );
  NAND2 U4472 ( .A(\mult_49/ab[1][6] ), .B(n317), .OUT(n2214) );
  NAND2 U4473 ( .A(n316), .B(n315), .OUT(n3740) );
  NAND2 U4474 ( .A(\mult_49/ab[2][6] ), .B(n5092), .OUT(n3739) );
  NAND2 U4475 ( .A(n2201), .B(n5650), .OUT(n2218) );
  NOR2 U4476 ( .A(n5650), .B(n2201), .OUT(n5651) );
  NOR2 U4477 ( .A(n5652), .B(n3754), .OUT(n2221) );
  NOR2 U4478 ( .A(n5653), .B(n2204), .OUT(n2220) );
  NOR2 U4479 ( .A(n2207), .B(n3771), .OUT(n5654) );
  NAND2 U4480 ( .A(n3771), .B(n2207), .OUT(n2223) );
  NOR2 U4481 ( .A(n2210), .B(n3792), .OUT(n5655) );
  NAND2 U4482 ( .A(n3792), .B(n2210), .OUT(n2226) );
  NAND2 U4483 ( .A(\mult_49/ab[0][6] ), .B(n334), .OUT(n2230) );
  NAND2 U4484 ( .A(\mult_49/ab[1][5] ), .B(n333), .OUT(n2229) );
  NAND2 U4485 ( .A(n332), .B(n331), .OUT(n3729) );
  NAND2 U4486 ( .A(\mult_49/ab[2][5] ), .B(n5093), .OUT(n3728) );
  NAND2 U4487 ( .A(n2213), .B(n5656), .OUT(n2233) );
  NOR2 U4488 ( .A(n5656), .B(n2213), .OUT(n5657) );
  NOR2 U4489 ( .A(n5658), .B(n3741), .OUT(n2236) );
  NOR2 U4490 ( .A(n5659), .B(n2216), .OUT(n2235) );
  NOR2 U4491 ( .A(n2219), .B(n3756), .OUT(n5660) );
  NAND2 U4492 ( .A(n3756), .B(n2219), .OUT(n2238) );
  NAND2 U4493 ( .A(n2222), .B(n5662), .OUT(n5661) );
  NOR2 U4494 ( .A(n5662), .B(n2222), .OUT(n2241) );
  NAND2 U4495 ( .A(n2225), .B(n5664), .OUT(n5663) );
  NOR2 U4496 ( .A(n5664), .B(n2225), .OUT(n2244) );
  NAND2 U4497 ( .A(\mult_49/ab[0][5] ), .B(n354), .OUT(n2248) );
  NAND2 U4498 ( .A(\mult_49/ab[1][4] ), .B(n353), .OUT(n2247) );
  NAND2 U4499 ( .A(n352), .B(n351), .OUT(n3720) );
  NAND2 U4500 ( .A(\mult_49/ab[2][4] ), .B(n5094), .OUT(n3719) );
  NAND2 U4501 ( .A(n2228), .B(n5665), .OUT(n2251) );
  NOR2 U4502 ( .A(n5665), .B(n2228), .OUT(n5666) );
  NOR2 U4503 ( .A(n5667), .B(n3730), .OUT(n2254) );
  NOR2 U4504 ( .A(n5668), .B(n2231), .OUT(n2253) );
  NOR2 U4505 ( .A(n2234), .B(n3743), .OUT(n5669) );
  NAND2 U4506 ( .A(n3743), .B(n2234), .OUT(n2256) );
  NAND2 U4507 ( .A(n2237), .B(n5671), .OUT(n5670) );
  NOR2 U4508 ( .A(n5671), .B(n2237), .OUT(n2259) );
  NOR2 U4509 ( .A(n2240), .B(n3775), .OUT(n5672) );
  NAND2 U4510 ( .A(n3775), .B(n2240), .OUT(n2262) );
  NOR2 U4511 ( .A(n2243), .B(n3796), .OUT(n5673) );
  NAND2 U4512 ( .A(n3796), .B(n2243), .OUT(n2265) );
  NAND2 U4513 ( .A(\mult_49/ab[0][4] ), .B(n378), .OUT(n2269) );
  NAND2 U4514 ( .A(\mult_49/ab[1][3] ), .B(n377), .OUT(n2268) );
  NAND2 U4515 ( .A(n376), .B(n375), .OUT(n3713) );
  NAND2 U4516 ( .A(\mult_49/ab[2][3] ), .B(n5095), .OUT(n3712) );
  NAND2 U4517 ( .A(n2246), .B(n5674), .OUT(n2272) );
  NOR2 U4518 ( .A(n5674), .B(n2246), .OUT(n5675) );
  NOR2 U4519 ( .A(n5676), .B(n3721), .OUT(n2275) );
  NOR2 U4520 ( .A(n5677), .B(n2249), .OUT(n2274) );
  NOR2 U4521 ( .A(n2252), .B(n3732), .OUT(n5678) );
  NAND2 U4522 ( .A(n3732), .B(n2252), .OUT(n2277) );
  NAND2 U4523 ( .A(n2255), .B(n5680), .OUT(n5679) );
  NOR2 U4524 ( .A(n5680), .B(n2255), .OUT(n2280) );
  NOR2 U4525 ( .A(n2258), .B(n3760), .OUT(n5681) );
  NAND2 U4526 ( .A(n3760), .B(n2258), .OUT(n2283) );
  NAND2 U4527 ( .A(n2261), .B(n5683), .OUT(n5682) );
  NOR2 U4528 ( .A(n5683), .B(n2261), .OUT(n2286) );
  NAND2 U4529 ( .A(n2264), .B(n5685), .OUT(n5684) );
  NOR2 U4530 ( .A(n5685), .B(n2264), .OUT(n2289) );
  NAND2 U4531 ( .A(\mult_49/ab[0][3] ), .B(n406), .OUT(n2293) );
  NAND2 U4532 ( .A(\mult_49/ab[1][2] ), .B(n405), .OUT(n2292) );
  NAND2 U4533 ( .A(n404), .B(n403), .OUT(n3708) );
  NAND2 U4534 ( .A(\mult_49/ab[2][2] ), .B(n5096), .OUT(n3707) );
  NAND2 U4535 ( .A(n2267), .B(n5686), .OUT(n2296) );
  NOR2 U4536 ( .A(n5686), .B(n2267), .OUT(n5687) );
  NOR2 U4537 ( .A(n5688), .B(n3714), .OUT(n2299) );
  NOR2 U4538 ( .A(n5689), .B(n2270), .OUT(n2298) );
  NOR2 U4539 ( .A(n2273), .B(n3723), .OUT(n5690) );
  NAND2 U4540 ( .A(n3723), .B(n2273), .OUT(n2301) );
  NAND2 U4541 ( .A(n2276), .B(n5692), .OUT(n5691) );
  NOR2 U4542 ( .A(n5692), .B(n2276), .OUT(n2304) );
  NOR2 U4543 ( .A(n2279), .B(n3747), .OUT(n5693) );
  NAND2 U4544 ( .A(n3747), .B(n2279), .OUT(n2307) );
  NAND2 U4545 ( .A(n2282), .B(n5695), .OUT(n5694) );
  NOR2 U4546 ( .A(n5695), .B(n2282), .OUT(n2310) );
  NOR2 U4547 ( .A(n2285), .B(n3779), .OUT(n5696) );
  NAND2 U4548 ( .A(n3779), .B(n2285), .OUT(n2313) );
  NOR2 U4549 ( .A(n2288), .B(n3800), .OUT(n2317) );
  NAND2 U4550 ( .A(n3800), .B(n2288), .OUT(n5697) );
  INV U4551 ( .IN(n2315), .OUT(n5519) );
  NAND2 U4552 ( .A(\mult_49/ab[0][2] ), .B(n438), .OUT(n2320) );
  NAND2 U4553 ( .A(\mult_49/ab[1][1] ), .B(n437), .OUT(n2319) );
  NAND2 U4554 ( .A(n436), .B(n435), .OUT(n3705) );
  NAND2 U4555 ( .A(\mult_49/ab[2][1] ), .B(n5097), .OUT(n3704) );
  NAND2 U4556 ( .A(n2291), .B(n5699), .OUT(n5698) );
  NOR2 U4557 ( .A(n5699), .B(n2291), .OUT(n2322) );
  NOR2 U4558 ( .A(n5700), .B(n3709), .OUT(n2326) );
  NOR2 U4559 ( .A(n5701), .B(n2294), .OUT(n2325) );
  NOR2 U4560 ( .A(n2297), .B(n3716), .OUT(n2329) );
  NAND2 U4561 ( .A(n3716), .B(n2297), .OUT(n5702) );
  INV U4562 ( .IN(n2327), .OUT(n5147) );
  NAND2 U4563 ( .A(n2300), .B(n5704), .OUT(n5703) );
  NOR2 U4564 ( .A(n5704), .B(n2300), .OUT(n2331) );
  NOR2 U4565 ( .A(n2303), .B(n3736), .OUT(n2335) );
  NAND2 U4566 ( .A(n3736), .B(n2303), .OUT(n5705) );
  INV U4567 ( .IN(n2333), .OUT(n5150) );
  NAND2 U4568 ( .A(n2306), .B(n5707), .OUT(n5706) );
  NOR2 U4569 ( .A(n5707), .B(n2306), .OUT(n2337) );
  NOR2 U4570 ( .A(n2309), .B(n3764), .OUT(n2341) );
  NAND2 U4571 ( .A(n3764), .B(n2309), .OUT(n5708) );
  INV U4572 ( .IN(n2339), .OUT(n5153) );
  NAND2 U4573 ( .A(n2312), .B(n5710), .OUT(n5709) );
  NOR2 U4574 ( .A(n5710), .B(n2312), .OUT(n2343) );
  NAND2 U4575 ( .A(\mult_49/ab[10][0] ), .B(n503), .OUT(n509) );
  NAND2 U4576 ( .A(n5154), .B(n506), .OUT(n3805) );
  NOR2 U4577 ( .A(n2342), .B(n3804), .OUT(n5711) );
  NAND2 U4578 ( .A(n3804), .B(n2342), .OUT(n2345) );
  NAND2 U4579 ( .A(\mult_49/ab[9][0] ), .B(n499), .OUT(n504) );
  NAND2 U4580 ( .A(n5152), .B(n502), .OUT(n3807) );
  NAND2 U4581 ( .A(\mult_49/ab[8][0] ), .B(n495), .OUT(n500) );
  NAND2 U4582 ( .A(n5151), .B(n498), .OUT(n3809) );
  NOR2 U4583 ( .A(n2336), .B(n3808), .OUT(n5712) );
  NAND2 U4584 ( .A(n3808), .B(n2336), .OUT(n2347) );
  NAND2 U4585 ( .A(\mult_49/ab[7][0] ), .B(n491), .OUT(n496) );
  NAND2 U4586 ( .A(n5149), .B(n494), .OUT(n3811) );
  NAND2 U4587 ( .A(\mult_49/ab[6][0] ), .B(n487), .OUT(n492) );
  NAND2 U4588 ( .A(n5148), .B(n490), .OUT(n3813) );
  NOR2 U4589 ( .A(n2330), .B(n3812), .OUT(n5713) );
  NAND2 U4590 ( .A(n3812), .B(n2330), .OUT(n2349) );
  NAND2 U4591 ( .A(\mult_49/ab[5][0] ), .B(n483), .OUT(n488) );
  NAND2 U4592 ( .A(n5146), .B(n486), .OUT(n3815) );
  NAND2 U4593 ( .A(\mult_49/ab[4][0] ), .B(n479), .OUT(n484) );
  NAND2 U4594 ( .A(n5145), .B(n482), .OUT(n3817) );
  NOR2 U4595 ( .A(n2324), .B(n3816), .OUT(n5714) );
  NAND2 U4596 ( .A(n3816), .B(n2324), .OUT(n2351) );
  NOR2 U4597 ( .A(n5715), .B(\mult_49/ab[30][1] ), .OUT(n4729) );
  NOR2 U4598 ( .A(n5716), .B(\mult_49/ab[29][2] ), .OUT(n4728) );
  NAND2 U4599 ( .A(\mult_49/ab[31][0] ), .B(n4727), .OUT(n4732) );
  NOR2 U4600 ( .A(n4727), .B(\mult_49/ab[31][0] ), .OUT(n5717) );
  NAND2 U4601 ( .A(\mult_49/ab[0][12] ), .B(n551), .OUT(n2355) );
  NAND2 U4602 ( .A(\mult_49/ab[1][11] ), .B(n552), .OUT(n2354) );
  NAND2 U4603 ( .A(n514), .B(n517), .OUT(n3820) );
  NAND2 U4604 ( .A(\mult_49/ab[2][10] ), .B(n5088), .OUT(n3819) );
  NAND2 U4605 ( .A(n2353), .B(n5718), .OUT(n2358) );
  NOR2 U4606 ( .A(n5718), .B(n2353), .OUT(n5719) );
  NOR2 U4607 ( .A(n5720), .B(n3821), .OUT(n2361) );
  NOR2 U4608 ( .A(n5721), .B(n2356), .OUT(n2360) );
  NOR2 U4609 ( .A(n2359), .B(n3823), .OUT(n5722) );
  NAND2 U4610 ( .A(n3823), .B(n2359), .OUT(n2363) );
  NAND2 U4611 ( .A(n2362), .B(n5724), .OUT(n5723) );
  NOR2 U4612 ( .A(n5724), .B(n2362), .OUT(n2366) );
  NOR2 U4613 ( .A(n2365), .B(n3827), .OUT(n5725) );
  NAND2 U4614 ( .A(n3827), .B(n2365), .OUT(n2369) );
  NAND2 U4615 ( .A(n2368), .B(n5727), .OUT(n5726) );
  NOR2 U4616 ( .A(n5727), .B(n2368), .OUT(n2372) );
  NOR2 U4617 ( .A(n2371), .B(n3831), .OUT(n5728) );
  NAND2 U4618 ( .A(n3831), .B(n2371), .OUT(n2375) );
  NAND2 U4619 ( .A(n2374), .B(n5730), .OUT(n5729) );
  NOR2 U4620 ( .A(n5730), .B(n2374), .OUT(n2378) );
  NAND2 U4621 ( .A(\mult_49/ab[0][13] ), .B(n591), .OUT(n2382) );
  NAND2 U4622 ( .A(\mult_49/ab[1][12] ), .B(n592), .OUT(n2381) );
  NAND2 U4623 ( .A(n550), .B(n553), .OUT(n3837) );
  NAND2 U4624 ( .A(\mult_49/ab[2][11] ), .B(n5087), .OUT(n3836) );
  NAND2 U4625 ( .A(n2380), .B(n5731), .OUT(n2385) );
  NOR2 U4626 ( .A(n5731), .B(n2380), .OUT(n5732) );
  NOR2 U4627 ( .A(n5733), .B(n3838), .OUT(n2388) );
  NOR2 U4628 ( .A(n5734), .B(n2383), .OUT(n2387) );
  NOR2 U4629 ( .A(n2386), .B(n3840), .OUT(n5735) );
  NAND2 U4630 ( .A(n3840), .B(n2386), .OUT(n2390) );
  NAND2 U4631 ( .A(n2389), .B(n5737), .OUT(n5736) );
  NOR2 U4632 ( .A(n5737), .B(n2389), .OUT(n2393) );
  NOR2 U4633 ( .A(n2392), .B(n3844), .OUT(n5738) );
  NAND2 U4634 ( .A(n3844), .B(n2392), .OUT(n2396) );
  NAND2 U4635 ( .A(n2395), .B(n5740), .OUT(n5739) );
  NOR2 U4636 ( .A(n5740), .B(n2395), .OUT(n2399) );
  NOR2 U4637 ( .A(n2398), .B(n3848), .OUT(n5741) );
  NAND2 U4638 ( .A(n3848), .B(n2398), .OUT(n2402) );
  NAND2 U4639 ( .A(n2401), .B(n5743), .OUT(n5742) );
  NOR2 U4640 ( .A(n5743), .B(n2401), .OUT(n2405) );
  NOR2 U4641 ( .A(n2404), .B(n3852), .OUT(n5744) );
  NAND2 U4642 ( .A(n3852), .B(n2404), .OUT(n2408) );
  NAND2 U4643 ( .A(\mult_49/ab[0][14] ), .B(n635), .OUT(n2412) );
  NAND2 U4644 ( .A(\mult_49/ab[1][13] ), .B(n636), .OUT(n2411) );
  NAND2 U4645 ( .A(n590), .B(n593), .OUT(n3856) );
  NAND2 U4646 ( .A(\mult_49/ab[2][12] ), .B(n5086), .OUT(n3855) );
  NAND2 U4647 ( .A(n2410), .B(n5745), .OUT(n2415) );
  NOR2 U4648 ( .A(n5745), .B(n2410), .OUT(n5746) );
  NOR2 U4649 ( .A(n5747), .B(n3857), .OUT(n2418) );
  NOR2 U4650 ( .A(n5748), .B(n2413), .OUT(n2417) );
  NOR2 U4651 ( .A(n2416), .B(n3859), .OUT(n5749) );
  NAND2 U4652 ( .A(n3859), .B(n2416), .OUT(n2420) );
  NAND2 U4653 ( .A(n2419), .B(n5751), .OUT(n5750) );
  NOR2 U4654 ( .A(n5751), .B(n2419), .OUT(n2423) );
  NOR2 U4655 ( .A(n2422), .B(n3863), .OUT(n5752) );
  NAND2 U4656 ( .A(n3863), .B(n2422), .OUT(n2426) );
  NAND2 U4657 ( .A(n2425), .B(n5754), .OUT(n5753) );
  NOR2 U4658 ( .A(n5754), .B(n2425), .OUT(n2429) );
  NOR2 U4659 ( .A(n2428), .B(n3867), .OUT(n5755) );
  NAND2 U4660 ( .A(n3867), .B(n2428), .OUT(n2432) );
  NAND2 U4661 ( .A(n2431), .B(n5757), .OUT(n5756) );
  NOR2 U4662 ( .A(n5757), .B(n2431), .OUT(n2435) );
  NOR2 U4663 ( .A(n2434), .B(n3871), .OUT(n5758) );
  NAND2 U4664 ( .A(n3871), .B(n2434), .OUT(n2438) );
  NAND2 U4665 ( .A(n2437), .B(n5760), .OUT(n5759) );
  NOR2 U4666 ( .A(n5760), .B(n2437), .OUT(n2441) );
  NAND2 U4667 ( .A(\mult_49/ab[0][15] ), .B(n683), .OUT(n2445) );
  NAND2 U4668 ( .A(\mult_49/ab[1][14] ), .B(n684), .OUT(n2444) );
  NAND2 U4669 ( .A(n634), .B(n637), .OUT(n3877) );
  NAND2 U4670 ( .A(\mult_49/ab[2][13] ), .B(n5085), .OUT(n3876) );
  NAND2 U4671 ( .A(n2443), .B(n5761), .OUT(n2448) );
  NOR2 U4672 ( .A(n5761), .B(n2443), .OUT(n5762) );
  NOR2 U4673 ( .A(n5763), .B(n3878), .OUT(n2451) );
  NOR2 U4674 ( .A(n5764), .B(n2446), .OUT(n2450) );
  NOR2 U4675 ( .A(n2449), .B(n3880), .OUT(n5765) );
  NAND2 U4676 ( .A(n3880), .B(n2449), .OUT(n2453) );
  NAND2 U4677 ( .A(n2452), .B(n5767), .OUT(n5766) );
  NOR2 U4678 ( .A(n5767), .B(n2452), .OUT(n2456) );
  NOR2 U4679 ( .A(n2455), .B(n3884), .OUT(n5768) );
  NAND2 U4680 ( .A(n3884), .B(n2455), .OUT(n2459) );
  NAND2 U4681 ( .A(n2458), .B(n5770), .OUT(n5769) );
  NOR2 U4682 ( .A(n5770), .B(n2458), .OUT(n2462) );
  NOR2 U4683 ( .A(n2461), .B(n3888), .OUT(n5771) );
  NAND2 U4684 ( .A(n3888), .B(n2461), .OUT(n2465) );
  NAND2 U4685 ( .A(n2464), .B(n5773), .OUT(n5772) );
  NOR2 U4686 ( .A(n5773), .B(n2464), .OUT(n2468) );
  NOR2 U4687 ( .A(n2467), .B(n3892), .OUT(n5774) );
  NAND2 U4688 ( .A(n3892), .B(n2467), .OUT(n2471) );
  NAND2 U4689 ( .A(n2470), .B(n5776), .OUT(n5775) );
  NOR2 U4690 ( .A(n5776), .B(n2470), .OUT(n2474) );
  NOR2 U4691 ( .A(n2473), .B(n3896), .OUT(n5777) );
  NAND2 U4692 ( .A(n3896), .B(n2473), .OUT(n2477) );
  NAND2 U4693 ( .A(\mult_49/ab[0][16] ), .B(n735), .OUT(n2481) );
  NAND2 U4694 ( .A(\mult_49/ab[1][15] ), .B(n736), .OUT(n2480) );
  NAND2 U4695 ( .A(n682), .B(n685), .OUT(n3900) );
  NAND2 U4696 ( .A(\mult_49/ab[2][14] ), .B(n5084), .OUT(n3899) );
  NAND2 U4697 ( .A(n2479), .B(n5778), .OUT(n2484) );
  NOR2 U4698 ( .A(n5778), .B(n2479), .OUT(n5779) );
  NOR2 U4699 ( .A(n5780), .B(n3901), .OUT(n2487) );
  NOR2 U4700 ( .A(n5781), .B(n2482), .OUT(n2486) );
  NOR2 U4701 ( .A(n2485), .B(n3903), .OUT(n5782) );
  NAND2 U4702 ( .A(n3903), .B(n2485), .OUT(n2489) );
  NAND2 U4703 ( .A(n2488), .B(n5784), .OUT(n5783) );
  NOR2 U4704 ( .A(n5784), .B(n2488), .OUT(n2492) );
  NOR2 U4705 ( .A(n2491), .B(n3907), .OUT(n5785) );
  NAND2 U4706 ( .A(n3907), .B(n2491), .OUT(n2495) );
  NAND2 U4707 ( .A(n2494), .B(n5787), .OUT(n5786) );
  NOR2 U4708 ( .A(n5787), .B(n2494), .OUT(n2498) );
  NOR2 U4709 ( .A(n2497), .B(n3911), .OUT(n5788) );
  NAND2 U4710 ( .A(n3911), .B(n2497), .OUT(n2501) );
  NAND2 U4711 ( .A(n2500), .B(n5790), .OUT(n5789) );
  NOR2 U4712 ( .A(n5790), .B(n2500), .OUT(n2504) );
  NOR2 U4713 ( .A(n2503), .B(n3915), .OUT(n5791) );
  NAND2 U4714 ( .A(n3915), .B(n2503), .OUT(n2507) );
  NAND2 U4715 ( .A(n2506), .B(n5793), .OUT(n5792) );
  NOR2 U4716 ( .A(n5793), .B(n2506), .OUT(n2510) );
  NOR2 U4717 ( .A(n2509), .B(n3919), .OUT(n5794) );
  NAND2 U4718 ( .A(n3919), .B(n2509), .OUT(n2513) );
  NAND2 U4719 ( .A(n2512), .B(n5796), .OUT(n5795) );
  NOR2 U4720 ( .A(n5796), .B(n2512), .OUT(n2516) );
  NAND2 U4721 ( .A(\mult_49/ab[0][17] ), .B(n791), .OUT(n2520) );
  NAND2 U4722 ( .A(\mult_49/ab[1][16] ), .B(n792), .OUT(n2519) );
  NAND2 U4723 ( .A(n734), .B(n737), .OUT(n3925) );
  NAND2 U4724 ( .A(\mult_49/ab[2][15] ), .B(n5083), .OUT(n3924) );
  NAND2 U4725 ( .A(n2518), .B(n5797), .OUT(n2523) );
  NOR2 U4726 ( .A(n5797), .B(n2518), .OUT(n5798) );
  NOR2 U4727 ( .A(n5799), .B(n3926), .OUT(n2526) );
  NOR2 U4728 ( .A(n5800), .B(n2521), .OUT(n2525) );
  NOR2 U4729 ( .A(n2524), .B(n3928), .OUT(n5801) );
  NAND2 U4730 ( .A(n3928), .B(n2524), .OUT(n2528) );
  NAND2 U4731 ( .A(n2527), .B(n5803), .OUT(n5802) );
  NOR2 U4732 ( .A(n5803), .B(n2527), .OUT(n2531) );
  NOR2 U4733 ( .A(n2530), .B(n3932), .OUT(n5804) );
  NAND2 U4734 ( .A(n3932), .B(n2530), .OUT(n2534) );
  NAND2 U4735 ( .A(n2533), .B(n5806), .OUT(n5805) );
  NOR2 U4736 ( .A(n5806), .B(n2533), .OUT(n2537) );
  NOR2 U4737 ( .A(n2536), .B(n3936), .OUT(n5807) );
  NAND2 U4738 ( .A(n3936), .B(n2536), .OUT(n2540) );
  NAND2 U4739 ( .A(n2539), .B(n5809), .OUT(n5808) );
  NOR2 U4740 ( .A(n5809), .B(n2539), .OUT(n2543) );
  NOR2 U4741 ( .A(n2542), .B(n3940), .OUT(n5810) );
  NAND2 U4742 ( .A(n3940), .B(n2542), .OUT(n2546) );
  NAND2 U4743 ( .A(n2545), .B(n5812), .OUT(n5811) );
  NOR2 U4744 ( .A(n5812), .B(n2545), .OUT(n2549) );
  NOR2 U4745 ( .A(n2548), .B(n3944), .OUT(n5813) );
  NAND2 U4746 ( .A(n3944), .B(n2548), .OUT(n2552) );
  NAND2 U4747 ( .A(n2551), .B(n5815), .OUT(n5814) );
  NOR2 U4748 ( .A(n5815), .B(n2551), .OUT(n2555) );
  NOR2 U4749 ( .A(n2554), .B(n3948), .OUT(n5816) );
  NAND2 U4750 ( .A(n3948), .B(n2554), .OUT(n2558) );
  NAND2 U4751 ( .A(\mult_49/ab[0][18] ), .B(n851), .OUT(n2562) );
  NAND2 U4752 ( .A(\mult_49/ab[1][17] ), .B(n852), .OUT(n2561) );
  NAND2 U4753 ( .A(n790), .B(n793), .OUT(n3952) );
  NAND2 U4754 ( .A(\mult_49/ab[2][16] ), .B(n5082), .OUT(n3951) );
  NAND2 U4755 ( .A(n2560), .B(n5817), .OUT(n2565) );
  NOR2 U4756 ( .A(n5817), .B(n2560), .OUT(n5818) );
  NOR2 U4757 ( .A(n5819), .B(n3953), .OUT(n2568) );
  NOR2 U4758 ( .A(n5820), .B(n2563), .OUT(n2567) );
  NOR2 U4759 ( .A(n2566), .B(n3955), .OUT(n5821) );
  NAND2 U4760 ( .A(n3955), .B(n2566), .OUT(n2570) );
  NAND2 U4761 ( .A(n2569), .B(n5823), .OUT(n5822) );
  NOR2 U4762 ( .A(n5823), .B(n2569), .OUT(n2573) );
  NOR2 U4763 ( .A(n2572), .B(n3959), .OUT(n5824) );
  NAND2 U4764 ( .A(n3959), .B(n2572), .OUT(n2576) );
  NAND2 U4765 ( .A(n2575), .B(n5826), .OUT(n5825) );
  NOR2 U4766 ( .A(n5826), .B(n2575), .OUT(n2579) );
  NOR2 U4767 ( .A(n2578), .B(n3963), .OUT(n5827) );
  NAND2 U4768 ( .A(n3963), .B(n2578), .OUT(n2582) );
  NAND2 U4769 ( .A(n2581), .B(n5829), .OUT(n5828) );
  NOR2 U4770 ( .A(n5829), .B(n2581), .OUT(n2585) );
  NOR2 U4771 ( .A(n2584), .B(n3967), .OUT(n5830) );
  NAND2 U4772 ( .A(n3967), .B(n2584), .OUT(n2588) );
  NAND2 U4773 ( .A(n2587), .B(n5832), .OUT(n5831) );
  NOR2 U4774 ( .A(n5832), .B(n2587), .OUT(n2591) );
  NOR2 U4775 ( .A(n2590), .B(n3971), .OUT(n5833) );
  NAND2 U4776 ( .A(n3971), .B(n2590), .OUT(n2594) );
  NAND2 U4777 ( .A(n2593), .B(n5835), .OUT(n5834) );
  NOR2 U4778 ( .A(n5835), .B(n2593), .OUT(n2597) );
  NOR2 U4779 ( .A(n2596), .B(n3975), .OUT(n5836) );
  NAND2 U4780 ( .A(n3975), .B(n2596), .OUT(n2600) );
  NAND2 U4781 ( .A(n2599), .B(n5838), .OUT(n5837) );
  NOR2 U4782 ( .A(n5838), .B(n2599), .OUT(n2603) );
  NAND2 U4783 ( .A(\mult_49/ab[0][19] ), .B(n915), .OUT(n2607) );
  NAND2 U4784 ( .A(\mult_49/ab[1][18] ), .B(n916), .OUT(n2606) );
  NAND2 U4785 ( .A(n850), .B(n853), .OUT(n3981) );
  NAND2 U4786 ( .A(\mult_49/ab[2][17] ), .B(n5081), .OUT(n3980) );
  NAND2 U4787 ( .A(n2605), .B(n5839), .OUT(n2610) );
  NOR2 U4788 ( .A(n5839), .B(n2605), .OUT(n5840) );
  NOR2 U4789 ( .A(n5841), .B(n3982), .OUT(n2613) );
  NOR2 U4790 ( .A(n5842), .B(n2608), .OUT(n2612) );
  NOR2 U4791 ( .A(n2611), .B(n3984), .OUT(n5843) );
  NAND2 U4792 ( .A(n3984), .B(n2611), .OUT(n2615) );
  NAND2 U4793 ( .A(n2614), .B(n5845), .OUT(n5844) );
  NOR2 U4794 ( .A(n5845), .B(n2614), .OUT(n2618) );
  NOR2 U4795 ( .A(n2617), .B(n3988), .OUT(n5846) );
  NAND2 U4796 ( .A(n3988), .B(n2617), .OUT(n2621) );
  NAND2 U4797 ( .A(n2620), .B(n5848), .OUT(n5847) );
  NOR2 U4798 ( .A(n5848), .B(n2620), .OUT(n2624) );
  NOR2 U4799 ( .A(n2623), .B(n3992), .OUT(n5849) );
  NAND2 U4800 ( .A(n3992), .B(n2623), .OUT(n2627) );
  NAND2 U4801 ( .A(n2626), .B(n5851), .OUT(n5850) );
  NOR2 U4802 ( .A(n5851), .B(n2626), .OUT(n2630) );
  NOR2 U4803 ( .A(n2629), .B(n3996), .OUT(n5852) );
  NAND2 U4804 ( .A(n3996), .B(n2629), .OUT(n2633) );
  NAND2 U4805 ( .A(n2632), .B(n5854), .OUT(n5853) );
  NOR2 U4806 ( .A(n5854), .B(n2632), .OUT(n2636) );
  NOR2 U4807 ( .A(n2635), .B(n4000), .OUT(n5855) );
  NAND2 U4808 ( .A(n4000), .B(n2635), .OUT(n2639) );
  NAND2 U4809 ( .A(n2638), .B(n5857), .OUT(n5856) );
  NOR2 U4810 ( .A(n5857), .B(n2638), .OUT(n2642) );
  NOR2 U4811 ( .A(n2641), .B(n4004), .OUT(n5858) );
  NAND2 U4812 ( .A(n4004), .B(n2641), .OUT(n2645) );
  NAND2 U4813 ( .A(n2644), .B(n5860), .OUT(n5859) );
  NOR2 U4814 ( .A(n5860), .B(n2644), .OUT(n2648) );
  NOR2 U4815 ( .A(n2647), .B(n4008), .OUT(n5861) );
  NAND2 U4816 ( .A(n4008), .B(n2647), .OUT(n2651) );
  NAND2 U4817 ( .A(\mult_49/ab[0][20] ), .B(n983), .OUT(n2655) );
  NAND2 U4818 ( .A(\mult_49/ab[1][19] ), .B(n984), .OUT(n2654) );
  NAND2 U4819 ( .A(n914), .B(n917), .OUT(n4012) );
  NAND2 U4820 ( .A(\mult_49/ab[2][18] ), .B(n5080), .OUT(n4011) );
  NAND2 U4821 ( .A(n2653), .B(n5862), .OUT(n2658) );
  NOR2 U4822 ( .A(n5862), .B(n2653), .OUT(n5863) );
  NOR2 U4823 ( .A(n5864), .B(n4013), .OUT(n2661) );
  NOR2 U4824 ( .A(n5865), .B(n2656), .OUT(n2660) );
  NOR2 U4825 ( .A(n2659), .B(n4015), .OUT(n5866) );
  NAND2 U4826 ( .A(n4015), .B(n2659), .OUT(n2663) );
  NAND2 U4827 ( .A(n2662), .B(n5868), .OUT(n5867) );
  NOR2 U4828 ( .A(n5868), .B(n2662), .OUT(n2666) );
  NOR2 U4829 ( .A(n2665), .B(n4019), .OUT(n5869) );
  NAND2 U4830 ( .A(n4019), .B(n2665), .OUT(n2669) );
  NAND2 U4831 ( .A(n2668), .B(n5871), .OUT(n5870) );
  NOR2 U4832 ( .A(n5871), .B(n2668), .OUT(n2672) );
  NOR2 U4833 ( .A(n2671), .B(n4023), .OUT(n5872) );
  NAND2 U4834 ( .A(n4023), .B(n2671), .OUT(n2675) );
  NAND2 U4835 ( .A(n2674), .B(n5874), .OUT(n5873) );
  NOR2 U4836 ( .A(n5874), .B(n2674), .OUT(n2678) );
  NOR2 U4837 ( .A(n2677), .B(n4027), .OUT(n5875) );
  NAND2 U4838 ( .A(n4027), .B(n2677), .OUT(n2681) );
  NAND2 U4839 ( .A(n2680), .B(n5877), .OUT(n5876) );
  NOR2 U4840 ( .A(n5877), .B(n2680), .OUT(n2684) );
  NOR2 U4841 ( .A(n2683), .B(n4031), .OUT(n5878) );
  NAND2 U4842 ( .A(n4031), .B(n2683), .OUT(n2687) );
  NAND2 U4843 ( .A(n2686), .B(n5880), .OUT(n5879) );
  NOR2 U4844 ( .A(n5880), .B(n2686), .OUT(n2690) );
  NOR2 U4845 ( .A(n2689), .B(n4035), .OUT(n5881) );
  NAND2 U4846 ( .A(n4035), .B(n2689), .OUT(n2693) );
  NAND2 U4847 ( .A(n2692), .B(n5883), .OUT(n5882) );
  NOR2 U4848 ( .A(n5883), .B(n2692), .OUT(n2696) );
  NOR2 U4849 ( .A(n2695), .B(n4039), .OUT(n5884) );
  NAND2 U4850 ( .A(n4039), .B(n2695), .OUT(n2699) );
  NAND2 U4851 ( .A(n2698), .B(n5886), .OUT(n5885) );
  NOR2 U4852 ( .A(n5886), .B(n2698), .OUT(n2702) );
  NAND2 U4853 ( .A(\mult_49/ab[0][21] ), .B(n1055), .OUT(n2706) );
  NAND2 U4854 ( .A(\mult_49/ab[1][20] ), .B(n1056), .OUT(n2705) );
  NAND2 U4855 ( .A(n982), .B(n985), .OUT(n4045) );
  NAND2 U4856 ( .A(\mult_49/ab[2][19] ), .B(n5079), .OUT(n4044) );
  NAND2 U4857 ( .A(n2704), .B(n5887), .OUT(n2709) );
  NOR2 U4858 ( .A(n5887), .B(n2704), .OUT(n5888) );
  NOR2 U4859 ( .A(n5889), .B(n4046), .OUT(n2712) );
  NOR2 U4860 ( .A(n5890), .B(n2707), .OUT(n2711) );
  NOR2 U4861 ( .A(n2710), .B(n4048), .OUT(n5891) );
  NAND2 U4862 ( .A(n4048), .B(n2710), .OUT(n2714) );
  NAND2 U4863 ( .A(n2713), .B(n5893), .OUT(n5892) );
  NOR2 U4864 ( .A(n5893), .B(n2713), .OUT(n2717) );
  NOR2 U4865 ( .A(n2716), .B(n4052), .OUT(n5894) );
  NAND2 U4866 ( .A(n4052), .B(n2716), .OUT(n2720) );
  NAND2 U4867 ( .A(n2719), .B(n5896), .OUT(n5895) );
  NOR2 U4868 ( .A(n5896), .B(n2719), .OUT(n2723) );
  NOR2 U4869 ( .A(n2722), .B(n4056), .OUT(n5897) );
  NAND2 U4870 ( .A(n4056), .B(n2722), .OUT(n2726) );
  NAND2 U4871 ( .A(n2725), .B(n5899), .OUT(n5898) );
  NOR2 U4872 ( .A(n5899), .B(n2725), .OUT(n2729) );
  NOR2 U4873 ( .A(n2728), .B(n4060), .OUT(n5900) );
  NAND2 U4874 ( .A(n4060), .B(n2728), .OUT(n2732) );
  NAND2 U4875 ( .A(n2731), .B(n5902), .OUT(n5901) );
  NOR2 U4876 ( .A(n5902), .B(n2731), .OUT(n2735) );
  NOR2 U4877 ( .A(n2734), .B(n4064), .OUT(n5903) );
  NAND2 U4878 ( .A(n4064), .B(n2734), .OUT(n2738) );
  NAND2 U4879 ( .A(n2737), .B(n5905), .OUT(n5904) );
  NOR2 U4880 ( .A(n5905), .B(n2737), .OUT(n2741) );
  NOR2 U4881 ( .A(n2740), .B(n4068), .OUT(n5906) );
  NAND2 U4882 ( .A(n4068), .B(n2740), .OUT(n2744) );
  NAND2 U4883 ( .A(n2743), .B(n5908), .OUT(n5907) );
  NOR2 U4884 ( .A(n5908), .B(n2743), .OUT(n2747) );
  NOR2 U4885 ( .A(n2746), .B(n4072), .OUT(n5909) );
  NAND2 U4886 ( .A(n4072), .B(n2746), .OUT(n2750) );
  NAND2 U4887 ( .A(n2749), .B(n5911), .OUT(n5910) );
  NOR2 U4888 ( .A(n5911), .B(n2749), .OUT(n2753) );
  NOR2 U4889 ( .A(n2752), .B(n4076), .OUT(n5912) );
  NAND2 U4890 ( .A(n4076), .B(n2752), .OUT(n2756) );
  NAND2 U4891 ( .A(\mult_49/ab[0][22] ), .B(n1131), .OUT(n2760) );
  NAND2 U4892 ( .A(\mult_49/ab[1][21] ), .B(n1132), .OUT(n2759) );
  NAND2 U4893 ( .A(n1054), .B(n1057), .OUT(n4080) );
  NAND2 U4894 ( .A(\mult_49/ab[2][20] ), .B(n5078), .OUT(n4079) );
  NAND2 U4895 ( .A(n2758), .B(n5913), .OUT(n2763) );
  NOR2 U4896 ( .A(n5913), .B(n2758), .OUT(n5914) );
  NOR2 U4897 ( .A(n5915), .B(n4081), .OUT(n2766) );
  NOR2 U4898 ( .A(n5916), .B(n2761), .OUT(n2765) );
  NOR2 U4899 ( .A(n2764), .B(n4083), .OUT(n5917) );
  NAND2 U4900 ( .A(n4083), .B(n2764), .OUT(n2768) );
  NAND2 U4901 ( .A(n2767), .B(n5919), .OUT(n5918) );
  NOR2 U4902 ( .A(n5919), .B(n2767), .OUT(n2771) );
  NOR2 U4903 ( .A(n2770), .B(n4087), .OUT(n5920) );
  NAND2 U4904 ( .A(n4087), .B(n2770), .OUT(n2774) );
  NAND2 U4905 ( .A(n2773), .B(n5922), .OUT(n5921) );
  NOR2 U4906 ( .A(n5922), .B(n2773), .OUT(n2777) );
  NOR2 U4907 ( .A(n2776), .B(n4091), .OUT(n5923) );
  NAND2 U4908 ( .A(n4091), .B(n2776), .OUT(n2780) );
  NAND2 U4909 ( .A(n2779), .B(n5925), .OUT(n5924) );
  NOR2 U4910 ( .A(n5925), .B(n2779), .OUT(n2783) );
  NOR2 U4911 ( .A(n2782), .B(n4095), .OUT(n5926) );
  NAND2 U4912 ( .A(n4095), .B(n2782), .OUT(n2786) );
  NAND2 U4913 ( .A(n2785), .B(n5928), .OUT(n5927) );
  NOR2 U4914 ( .A(n5928), .B(n2785), .OUT(n2789) );
  NOR2 U4915 ( .A(n2788), .B(n4099), .OUT(n5929) );
  NAND2 U4916 ( .A(n4099), .B(n2788), .OUT(n2792) );
  NAND2 U4917 ( .A(n2791), .B(n5931), .OUT(n5930) );
  NOR2 U4918 ( .A(n5931), .B(n2791), .OUT(n2795) );
  NOR2 U4919 ( .A(n2794), .B(n4103), .OUT(n5932) );
  NAND2 U4920 ( .A(n4103), .B(n2794), .OUT(n2798) );
  NAND2 U4921 ( .A(n2797), .B(n5934), .OUT(n5933) );
  NOR2 U4922 ( .A(n5934), .B(n2797), .OUT(n2801) );
  NOR2 U4923 ( .A(n2800), .B(n4107), .OUT(n5935) );
  NAND2 U4924 ( .A(n4107), .B(n2800), .OUT(n2804) );
  NAND2 U4925 ( .A(n2803), .B(n5937), .OUT(n5936) );
  NOR2 U4926 ( .A(n5937), .B(n2803), .OUT(n2807) );
  NOR2 U4927 ( .A(n2806), .B(n4111), .OUT(n5938) );
  NAND2 U4928 ( .A(n4111), .B(n2806), .OUT(n2810) );
  NAND2 U4929 ( .A(n2809), .B(n5940), .OUT(n5939) );
  NOR2 U4930 ( .A(n5940), .B(n2809), .OUT(n2813) );
  NAND2 U4931 ( .A(\mult_49/ab[0][23] ), .B(n1211), .OUT(n2817) );
  NAND2 U4932 ( .A(\mult_49/ab[1][22] ), .B(n1212), .OUT(n2816) );
  NAND2 U4933 ( .A(n1130), .B(n1133), .OUT(n4117) );
  NAND2 U4934 ( .A(\mult_49/ab[2][21] ), .B(n5077), .OUT(n4116) );
  NAND2 U4935 ( .A(n2815), .B(n5941), .OUT(n2820) );
  NOR2 U4936 ( .A(n5941), .B(n2815), .OUT(n5942) );
  NOR2 U4937 ( .A(n5943), .B(n4118), .OUT(n2823) );
  NOR2 U4938 ( .A(n5944), .B(n2818), .OUT(n2822) );
  NOR2 U4939 ( .A(n2821), .B(n4120), .OUT(n5945) );
  NAND2 U4940 ( .A(n4120), .B(n2821), .OUT(n2825) );
  NAND2 U4941 ( .A(n2824), .B(n5947), .OUT(n5946) );
  NOR2 U4942 ( .A(n5947), .B(n2824), .OUT(n2828) );
  NOR2 U4943 ( .A(n2827), .B(n4124), .OUT(n5948) );
  NAND2 U4944 ( .A(n4124), .B(n2827), .OUT(n2831) );
  NAND2 U4945 ( .A(n2830), .B(n5950), .OUT(n5949) );
  NOR2 U4946 ( .A(n5950), .B(n2830), .OUT(n2834) );
  NOR2 U4947 ( .A(n2833), .B(n4128), .OUT(n5951) );
  NAND2 U4948 ( .A(n4128), .B(n2833), .OUT(n2837) );
  NAND2 U4949 ( .A(n2836), .B(n5953), .OUT(n5952) );
  NOR2 U4950 ( .A(n5953), .B(n2836), .OUT(n2840) );
  NOR2 U4951 ( .A(n2839), .B(n4132), .OUT(n5954) );
  NAND2 U4952 ( .A(n4132), .B(n2839), .OUT(n2843) );
  NAND2 U4953 ( .A(n2842), .B(n5956), .OUT(n5955) );
  NOR2 U4954 ( .A(n5956), .B(n2842), .OUT(n2846) );
  NOR2 U4955 ( .A(n2845), .B(n4136), .OUT(n5957) );
  NAND2 U4956 ( .A(n4136), .B(n2845), .OUT(n2849) );
  NAND2 U4957 ( .A(n2848), .B(n5959), .OUT(n5958) );
  NOR2 U4958 ( .A(n5959), .B(n2848), .OUT(n2852) );
  NOR2 U4959 ( .A(n2851), .B(n4140), .OUT(n5960) );
  NAND2 U4960 ( .A(n4140), .B(n2851), .OUT(n2855) );
  NAND2 U4961 ( .A(n2854), .B(n5962), .OUT(n5961) );
  NOR2 U4962 ( .A(n5962), .B(n2854), .OUT(n2858) );
  NOR2 U4963 ( .A(n2857), .B(n4144), .OUT(n5963) );
  NAND2 U4964 ( .A(n4144), .B(n2857), .OUT(n2861) );
  NAND2 U4965 ( .A(n2860), .B(n5965), .OUT(n5964) );
  NOR2 U4966 ( .A(n5965), .B(n2860), .OUT(n2864) );
  NOR2 U4967 ( .A(n2863), .B(n4148), .OUT(n5966) );
  NAND2 U4968 ( .A(n4148), .B(n2863), .OUT(n2867) );
  NAND2 U4969 ( .A(n2866), .B(n5968), .OUT(n5967) );
  NOR2 U4970 ( .A(n5968), .B(n2866), .OUT(n2870) );
  NOR2 U4971 ( .A(n2869), .B(n4152), .OUT(n5969) );
  NAND2 U4972 ( .A(n4152), .B(n2869), .OUT(n2873) );
  NAND2 U4973 ( .A(\mult_49/ab[0][24] ), .B(n1295), .OUT(n2877) );
  NAND2 U4974 ( .A(\mult_49/ab[1][23] ), .B(n1296), .OUT(n2876) );
  NAND2 U4975 ( .A(n1210), .B(n1213), .OUT(n4156) );
  NAND2 U4976 ( .A(\mult_49/ab[2][22] ), .B(n5076), .OUT(n4155) );
  NAND2 U4977 ( .A(n2875), .B(n5970), .OUT(n2880) );
  NOR2 U4978 ( .A(n5970), .B(n2875), .OUT(n5971) );
  NOR2 U4979 ( .A(n5972), .B(n4157), .OUT(n2883) );
  NOR2 U4980 ( .A(n5973), .B(n2878), .OUT(n2882) );
  NOR2 U4981 ( .A(n2881), .B(n4159), .OUT(n5974) );
  NAND2 U4982 ( .A(n4159), .B(n2881), .OUT(n2885) );
  NAND2 U4983 ( .A(n2884), .B(n5976), .OUT(n5975) );
  NOR2 U4984 ( .A(n5976), .B(n2884), .OUT(n2888) );
  NOR2 U4985 ( .A(n2887), .B(n4163), .OUT(n5977) );
  NAND2 U4986 ( .A(n4163), .B(n2887), .OUT(n2891) );
  NAND2 U4987 ( .A(n2890), .B(n5979), .OUT(n5978) );
  NOR2 U4988 ( .A(n5979), .B(n2890), .OUT(n2894) );
  NOR2 U4989 ( .A(n2893), .B(n4167), .OUT(n5980) );
  NAND2 U4990 ( .A(n4167), .B(n2893), .OUT(n2897) );
  NAND2 U4991 ( .A(n2896), .B(n5982), .OUT(n5981) );
  NOR2 U4992 ( .A(n5982), .B(n2896), .OUT(n2900) );
  NOR2 U4993 ( .A(n2899), .B(n4171), .OUT(n5983) );
  NAND2 U4994 ( .A(n4171), .B(n2899), .OUT(n2903) );
  NAND2 U4995 ( .A(n2902), .B(n5985), .OUT(n5984) );
  NOR2 U4996 ( .A(n5985), .B(n2902), .OUT(n2906) );
  NOR2 U4997 ( .A(n2905), .B(n4175), .OUT(n5986) );
  NAND2 U4998 ( .A(n4175), .B(n2905), .OUT(n2909) );
  NAND2 U4999 ( .A(n2908), .B(n5988), .OUT(n5987) );
  NOR2 U5000 ( .A(n5988), .B(n2908), .OUT(n2912) );
  NOR2 U5001 ( .A(n2911), .B(n4179), .OUT(n5989) );
  NAND2 U5002 ( .A(n4179), .B(n2911), .OUT(n2915) );
  NAND2 U5003 ( .A(n2914), .B(n5991), .OUT(n5990) );
  NOR2 U5004 ( .A(n5991), .B(n2914), .OUT(n2918) );
  NOR2 U5005 ( .A(n2917), .B(n4183), .OUT(n5992) );
  NAND2 U5006 ( .A(n4183), .B(n2917), .OUT(n2921) );
  NAND2 U5007 ( .A(n2920), .B(n5994), .OUT(n5993) );
  NOR2 U5008 ( .A(n5994), .B(n2920), .OUT(n2924) );
  NOR2 U5009 ( .A(n2923), .B(n4187), .OUT(n5995) );
  NAND2 U5010 ( .A(n4187), .B(n2923), .OUT(n2927) );
  NAND2 U5011 ( .A(n2926), .B(n5997), .OUT(n5996) );
  NOR2 U5012 ( .A(n5997), .B(n2926), .OUT(n2930) );
  NOR2 U5013 ( .A(n2929), .B(n4191), .OUT(n5998) );
  NAND2 U5014 ( .A(n4191), .B(n2929), .OUT(n2933) );
  NAND2 U5015 ( .A(n2932), .B(n6000), .OUT(n5999) );
  NOR2 U5016 ( .A(n6000), .B(n2932), .OUT(n2936) );
  NAND2 U5017 ( .A(\mult_49/ab[0][25] ), .B(n1383), .OUT(n2940) );
  NAND2 U5018 ( .A(\mult_49/ab[1][24] ), .B(n1384), .OUT(n2939) );
  NAND2 U5019 ( .A(n1294), .B(n1297), .OUT(n4197) );
  NAND2 U5020 ( .A(\mult_49/ab[2][23] ), .B(n5075), .OUT(n4196) );
  NAND2 U5021 ( .A(n2938), .B(n6001), .OUT(n2943) );
  NOR2 U5022 ( .A(n6001), .B(n2938), .OUT(n6002) );
  NOR2 U5023 ( .A(n6003), .B(n4198), .OUT(n2946) );
  NOR2 U5024 ( .A(n6004), .B(n2941), .OUT(n2945) );
  NOR2 U5025 ( .A(n2944), .B(n4200), .OUT(n6005) );
  NAND2 U5026 ( .A(n4200), .B(n2944), .OUT(n2948) );
  NAND2 U5027 ( .A(n2947), .B(n6007), .OUT(n6006) );
  NOR2 U5028 ( .A(n6007), .B(n2947), .OUT(n2951) );
  NOR2 U5029 ( .A(n2950), .B(n4204), .OUT(n6008) );
  NAND2 U5030 ( .A(n4204), .B(n2950), .OUT(n2954) );
  NAND2 U5031 ( .A(n2953), .B(n6010), .OUT(n6009) );
  NOR2 U5032 ( .A(n6010), .B(n2953), .OUT(n2957) );
  NOR2 U5033 ( .A(n2956), .B(n4208), .OUT(n6011) );
  NAND2 U5034 ( .A(n4208), .B(n2956), .OUT(n2960) );
  NAND2 U5035 ( .A(n2959), .B(n6013), .OUT(n6012) );
  NOR2 U5036 ( .A(n6013), .B(n2959), .OUT(n2963) );
  NOR2 U5037 ( .A(n2962), .B(n4212), .OUT(n6014) );
  NAND2 U5038 ( .A(n4212), .B(n2962), .OUT(n2966) );
  NAND2 U5039 ( .A(n2965), .B(n6016), .OUT(n6015) );
  NOR2 U5040 ( .A(n6016), .B(n2965), .OUT(n2969) );
  NOR2 U5041 ( .A(n2968), .B(n4216), .OUT(n6017) );
  NAND2 U5042 ( .A(n4216), .B(n2968), .OUT(n2972) );
  NAND2 U5043 ( .A(n2971), .B(n6019), .OUT(n6018) );
  NOR2 U5044 ( .A(n6019), .B(n2971), .OUT(n2975) );
  NOR2 U5045 ( .A(n2974), .B(n4220), .OUT(n6020) );
  NAND2 U5046 ( .A(n4220), .B(n2974), .OUT(n2978) );
  NAND2 U5047 ( .A(n2977), .B(n6022), .OUT(n6021) );
  NOR2 U5048 ( .A(n6022), .B(n2977), .OUT(n2981) );
  NOR2 U5049 ( .A(n2980), .B(n4224), .OUT(n6023) );
  NAND2 U5050 ( .A(n4224), .B(n2980), .OUT(n2984) );
  NAND2 U5051 ( .A(n2983), .B(n6025), .OUT(n6024) );
  NOR2 U5052 ( .A(n6025), .B(n2983), .OUT(n2987) );
  NOR2 U5053 ( .A(n2986), .B(n4228), .OUT(n6026) );
  NAND2 U5054 ( .A(n4228), .B(n2986), .OUT(n2990) );
  NAND2 U5055 ( .A(n2989), .B(n6028), .OUT(n6027) );
  NOR2 U5056 ( .A(n6028), .B(n2989), .OUT(n2993) );
  NOR2 U5057 ( .A(n2992), .B(n4232), .OUT(n6029) );
  NAND2 U5058 ( .A(n4232), .B(n2992), .OUT(n2996) );
  NAND2 U5059 ( .A(n2995), .B(n6031), .OUT(n6030) );
  NOR2 U5060 ( .A(n6031), .B(n2995), .OUT(n2999) );
  NOR2 U5061 ( .A(n2998), .B(n4236), .OUT(n6032) );
  NAND2 U5062 ( .A(n4236), .B(n2998), .OUT(n3002) );
  NAND2 U5063 ( .A(\mult_49/ab[0][26] ), .B(n1475), .OUT(n3006) );
  NAND2 U5064 ( .A(\mult_49/ab[1][25] ), .B(n1476), .OUT(n3005) );
  NAND2 U5065 ( .A(n1382), .B(n1385), .OUT(n4240) );
  NAND2 U5066 ( .A(\mult_49/ab[2][24] ), .B(n5074), .OUT(n4239) );
  NAND2 U5067 ( .A(n3004), .B(n6033), .OUT(n3009) );
  NOR2 U5068 ( .A(n6033), .B(n3004), .OUT(n6034) );
  NOR2 U5069 ( .A(n6035), .B(n4241), .OUT(n3012) );
  NOR2 U5070 ( .A(n6036), .B(n3007), .OUT(n3011) );
  NOR2 U5071 ( .A(n3010), .B(n4243), .OUT(n6037) );
  NAND2 U5072 ( .A(n4243), .B(n3010), .OUT(n3014) );
  NAND2 U5073 ( .A(n3013), .B(n6039), .OUT(n6038) );
  NOR2 U5074 ( .A(n6039), .B(n3013), .OUT(n3017) );
  NOR2 U5075 ( .A(n3016), .B(n4247), .OUT(n6040) );
  NAND2 U5076 ( .A(n4247), .B(n3016), .OUT(n3020) );
  NAND2 U5077 ( .A(n3019), .B(n6042), .OUT(n6041) );
  NOR2 U5078 ( .A(n6042), .B(n3019), .OUT(n3023) );
  NOR2 U5079 ( .A(n3022), .B(n4251), .OUT(n6043) );
  NAND2 U5080 ( .A(n4251), .B(n3022), .OUT(n3026) );
  NAND2 U5081 ( .A(n3025), .B(n6045), .OUT(n6044) );
  NOR2 U5082 ( .A(n6045), .B(n3025), .OUT(n3029) );
  NOR2 U5083 ( .A(n3028), .B(n4255), .OUT(n6046) );
  NAND2 U5084 ( .A(n4255), .B(n3028), .OUT(n3032) );
  NAND2 U5085 ( .A(n3031), .B(n6048), .OUT(n6047) );
  NOR2 U5086 ( .A(n6048), .B(n3031), .OUT(n3035) );
  NOR2 U5087 ( .A(n3034), .B(n4259), .OUT(n6049) );
  NAND2 U5088 ( .A(n4259), .B(n3034), .OUT(n3038) );
  NAND2 U5089 ( .A(n3037), .B(n6051), .OUT(n6050) );
  NOR2 U5090 ( .A(n6051), .B(n3037), .OUT(n3041) );
  NOR2 U5091 ( .A(n3040), .B(n4263), .OUT(n6052) );
  NAND2 U5092 ( .A(n4263), .B(n3040), .OUT(n3044) );
  NAND2 U5093 ( .A(n3043), .B(n6054), .OUT(n6053) );
  NOR2 U5094 ( .A(n6054), .B(n3043), .OUT(n3047) );
  NOR2 U5095 ( .A(n3046), .B(n4267), .OUT(n6055) );
  NAND2 U5096 ( .A(n4267), .B(n3046), .OUT(n3050) );
  NAND2 U5097 ( .A(n3049), .B(n6057), .OUT(n6056) );
  NOR2 U5098 ( .A(n6057), .B(n3049), .OUT(n3053) );
  NOR2 U5099 ( .A(n3052), .B(n4271), .OUT(n6058) );
  NAND2 U5100 ( .A(n4271), .B(n3052), .OUT(n3056) );
  NAND2 U5101 ( .A(n3055), .B(n6060), .OUT(n6059) );
  NOR2 U5102 ( .A(n6060), .B(n3055), .OUT(n3059) );
  NOR2 U5103 ( .A(n3058), .B(n4275), .OUT(n6061) );
  NAND2 U5104 ( .A(n4275), .B(n3058), .OUT(n3062) );
  NAND2 U5105 ( .A(n3061), .B(n6063), .OUT(n6062) );
  NOR2 U5106 ( .A(n6063), .B(n3061), .OUT(n3065) );
  NOR2 U5107 ( .A(n3064), .B(n4279), .OUT(n6064) );
  NAND2 U5108 ( .A(n4279), .B(n3064), .OUT(n3068) );
  NAND2 U5109 ( .A(n3067), .B(n6066), .OUT(n6065) );
  NOR2 U5110 ( .A(n6066), .B(n3067), .OUT(n3071) );
  NAND2 U5111 ( .A(\mult_49/ab[0][27] ), .B(n1571), .OUT(n3075) );
  NAND2 U5112 ( .A(\mult_49/ab[1][26] ), .B(n1572), .OUT(n3074) );
  NAND2 U5113 ( .A(n1474), .B(n1477), .OUT(n4285) );
  NAND2 U5114 ( .A(\mult_49/ab[2][25] ), .B(n5073), .OUT(n4284) );
  NAND2 U5115 ( .A(n3073), .B(n6067), .OUT(n3078) );
  NOR2 U5116 ( .A(n6067), .B(n3073), .OUT(n6068) );
  NOR2 U5117 ( .A(n6069), .B(n4286), .OUT(n3081) );
  NOR2 U5118 ( .A(n6070), .B(n3076), .OUT(n3080) );
  NOR2 U5119 ( .A(n3079), .B(n4288), .OUT(n6071) );
  NAND2 U5120 ( .A(n4288), .B(n3079), .OUT(n3083) );
  NAND2 U5121 ( .A(n3082), .B(n6073), .OUT(n6072) );
  NOR2 U5122 ( .A(n6073), .B(n3082), .OUT(n3086) );
  NOR2 U5123 ( .A(n3085), .B(n4292), .OUT(n6074) );
  NAND2 U5124 ( .A(n4292), .B(n3085), .OUT(n3089) );
  NAND2 U5125 ( .A(n3088), .B(n6076), .OUT(n6075) );
  NOR2 U5126 ( .A(n6076), .B(n3088), .OUT(n3092) );
  NOR2 U5127 ( .A(n3091), .B(n4296), .OUT(n6077) );
  NAND2 U5128 ( .A(n4296), .B(n3091), .OUT(n3095) );
  NAND2 U5129 ( .A(n3094), .B(n6079), .OUT(n6078) );
  NOR2 U5130 ( .A(n6079), .B(n3094), .OUT(n3098) );
  NOR2 U5131 ( .A(n3097), .B(n4300), .OUT(n6080) );
  NAND2 U5132 ( .A(n4300), .B(n3097), .OUT(n3101) );
  NAND2 U5133 ( .A(n3100), .B(n6082), .OUT(n6081) );
  NOR2 U5134 ( .A(n6082), .B(n3100), .OUT(n3104) );
  NOR2 U5135 ( .A(n3103), .B(n4304), .OUT(n6083) );
  NAND2 U5136 ( .A(n4304), .B(n3103), .OUT(n3107) );
  NAND2 U5137 ( .A(n3106), .B(n6085), .OUT(n6084) );
  NOR2 U5138 ( .A(n6085), .B(n3106), .OUT(n3110) );
  NOR2 U5139 ( .A(n3109), .B(n4308), .OUT(n6086) );
  NAND2 U5140 ( .A(n4308), .B(n3109), .OUT(n3113) );
  NAND2 U5141 ( .A(n3112), .B(n6088), .OUT(n6087) );
  NOR2 U5142 ( .A(n6088), .B(n3112), .OUT(n3116) );
  NOR2 U5143 ( .A(n3115), .B(n4312), .OUT(n6089) );
  NAND2 U5144 ( .A(n4312), .B(n3115), .OUT(n3119) );
  NAND2 U5145 ( .A(n3118), .B(n6091), .OUT(n6090) );
  NOR2 U5146 ( .A(n6091), .B(n3118), .OUT(n3122) );
  NOR2 U5147 ( .A(n3121), .B(n4316), .OUT(n6092) );
  NAND2 U5148 ( .A(n4316), .B(n3121), .OUT(n3125) );
  NAND2 U5149 ( .A(n3124), .B(n6094), .OUT(n6093) );
  NOR2 U5150 ( .A(n6094), .B(n3124), .OUT(n3128) );
  NOR2 U5151 ( .A(n3127), .B(n4320), .OUT(n6095) );
  NAND2 U5152 ( .A(n4320), .B(n3127), .OUT(n3131) );
  NAND2 U5153 ( .A(n3130), .B(n6097), .OUT(n6096) );
  NOR2 U5154 ( .A(n6097), .B(n3130), .OUT(n3134) );
  NOR2 U5155 ( .A(n3133), .B(n4324), .OUT(n6098) );
  NAND2 U5156 ( .A(n4324), .B(n3133), .OUT(n3137) );
  NAND2 U5157 ( .A(n3136), .B(n6100), .OUT(n6099) );
  NOR2 U5158 ( .A(n6100), .B(n3136), .OUT(n3140) );
  NOR2 U5159 ( .A(n3139), .B(n4328), .OUT(n6101) );
  NAND2 U5160 ( .A(n4328), .B(n3139), .OUT(n3143) );
  NAND2 U5161 ( .A(\mult_49/ab[0][28] ), .B(n1671), .OUT(n3147) );
  NAND2 U5162 ( .A(\mult_49/ab[1][27] ), .B(n1672), .OUT(n3146) );
  NAND2 U5163 ( .A(n1570), .B(n1573), .OUT(n4332) );
  NAND2 U5164 ( .A(\mult_49/ab[2][26] ), .B(n5072), .OUT(n4331) );
  NAND2 U5165 ( .A(n3145), .B(n6102), .OUT(n3150) );
  NOR2 U5166 ( .A(n6102), .B(n3145), .OUT(n6103) );
  NOR2 U5167 ( .A(n6104), .B(n4333), .OUT(n3153) );
  NOR2 U5168 ( .A(n6105), .B(n3148), .OUT(n3152) );
  NOR2 U5169 ( .A(n3151), .B(n4335), .OUT(n6106) );
  NAND2 U5170 ( .A(n4335), .B(n3151), .OUT(n3155) );
  NAND2 U5171 ( .A(n3154), .B(n6108), .OUT(n6107) );
  NOR2 U5172 ( .A(n6108), .B(n3154), .OUT(n3158) );
  NOR2 U5173 ( .A(n3157), .B(n4339), .OUT(n6109) );
  NAND2 U5174 ( .A(n4339), .B(n3157), .OUT(n3161) );
  NAND2 U5175 ( .A(n3160), .B(n6111), .OUT(n6110) );
  NOR2 U5176 ( .A(n6111), .B(n3160), .OUT(n3164) );
  NOR2 U5177 ( .A(n3163), .B(n4343), .OUT(n6112) );
  NAND2 U5178 ( .A(n4343), .B(n3163), .OUT(n3167) );
  NAND2 U5179 ( .A(n3166), .B(n6114), .OUT(n6113) );
  NOR2 U5180 ( .A(n6114), .B(n3166), .OUT(n3170) );
  NOR2 U5181 ( .A(n3169), .B(n4347), .OUT(n6115) );
  NAND2 U5182 ( .A(n4347), .B(n3169), .OUT(n3173) );
  NAND2 U5183 ( .A(n3172), .B(n6117), .OUT(n6116) );
  NOR2 U5184 ( .A(n6117), .B(n3172), .OUT(n3176) );
  NOR2 U5185 ( .A(n3175), .B(n4351), .OUT(n6118) );
  NAND2 U5186 ( .A(n4351), .B(n3175), .OUT(n3179) );
  NAND2 U5187 ( .A(n3178), .B(n6120), .OUT(n6119) );
  NOR2 U5188 ( .A(n6120), .B(n3178), .OUT(n3182) );
  NOR2 U5189 ( .A(n3181), .B(n4355), .OUT(n6121) );
  NAND2 U5190 ( .A(n4355), .B(n3181), .OUT(n3185) );
  NAND2 U5191 ( .A(n3184), .B(n6123), .OUT(n6122) );
  NOR2 U5192 ( .A(n6123), .B(n3184), .OUT(n3188) );
  NOR2 U5193 ( .A(n3187), .B(n4359), .OUT(n6124) );
  NAND2 U5194 ( .A(n4359), .B(n3187), .OUT(n3191) );
  NAND2 U5195 ( .A(n3190), .B(n6126), .OUT(n6125) );
  NOR2 U5196 ( .A(n6126), .B(n3190), .OUT(n3194) );
  NOR2 U5197 ( .A(n3193), .B(n4363), .OUT(n6127) );
  NAND2 U5198 ( .A(n4363), .B(n3193), .OUT(n3197) );
  NAND2 U5199 ( .A(n3196), .B(n6129), .OUT(n6128) );
  NOR2 U5200 ( .A(n6129), .B(n3196), .OUT(n3200) );
  NOR2 U5201 ( .A(n3199), .B(n4367), .OUT(n6130) );
  NAND2 U5202 ( .A(n4367), .B(n3199), .OUT(n3203) );
  NAND2 U5203 ( .A(n3202), .B(n6132), .OUT(n6131) );
  NOR2 U5204 ( .A(n6132), .B(n3202), .OUT(n3206) );
  NOR2 U5205 ( .A(n3205), .B(n4371), .OUT(n6133) );
  NAND2 U5206 ( .A(n4371), .B(n3205), .OUT(n3209) );
  NAND2 U5207 ( .A(n3208), .B(n6135), .OUT(n6134) );
  NOR2 U5208 ( .A(n6135), .B(n3208), .OUT(n3212) );
  NOR2 U5209 ( .A(n3211), .B(n4375), .OUT(n6136) );
  NAND2 U5210 ( .A(n4375), .B(n3211), .OUT(n3215) );
  NAND2 U5211 ( .A(n3214), .B(n6138), .OUT(n6137) );
  NOR2 U5212 ( .A(n6138), .B(n3214), .OUT(n3218) );
  NAND2 U5213 ( .A(\mult_49/ab[0][29] ), .B(n1775), .OUT(n3222) );
  NAND2 U5214 ( .A(\mult_49/ab[1][28] ), .B(n1776), .OUT(n3221) );
  NAND2 U5215 ( .A(n1670), .B(n1673), .OUT(n4381) );
  NAND2 U5216 ( .A(\mult_49/ab[2][27] ), .B(n5071), .OUT(n4380) );
  NAND2 U5217 ( .A(n3220), .B(n6139), .OUT(n3225) );
  NOR2 U5218 ( .A(n6139), .B(n3220), .OUT(n6140) );
  NOR2 U5219 ( .A(n6141), .B(n4382), .OUT(n3228) );
  NOR2 U5220 ( .A(n6142), .B(n3223), .OUT(n3227) );
  NOR2 U5221 ( .A(n3226), .B(n4384), .OUT(n6143) );
  NAND2 U5222 ( .A(n4384), .B(n3226), .OUT(n3230) );
  NAND2 U5223 ( .A(n3229), .B(n6145), .OUT(n6144) );
  NOR2 U5224 ( .A(n6145), .B(n3229), .OUT(n3233) );
  NOR2 U5225 ( .A(n3232), .B(n4388), .OUT(n6146) );
  NAND2 U5226 ( .A(n4388), .B(n3232), .OUT(n3236) );
  NAND2 U5227 ( .A(n3235), .B(n6148), .OUT(n6147) );
  NOR2 U5228 ( .A(n6148), .B(n3235), .OUT(n3239) );
  NOR2 U5229 ( .A(n3238), .B(n4392), .OUT(n6149) );
  NAND2 U5230 ( .A(n4392), .B(n3238), .OUT(n3242) );
  NAND2 U5231 ( .A(n3241), .B(n6151), .OUT(n6150) );
  NOR2 U5232 ( .A(n6151), .B(n3241), .OUT(n3245) );
  NOR2 U5233 ( .A(n3244), .B(n4396), .OUT(n6152) );
  NAND2 U5234 ( .A(n4396), .B(n3244), .OUT(n3248) );
  NAND2 U5235 ( .A(n3247), .B(n6154), .OUT(n6153) );
  NOR2 U5236 ( .A(n6154), .B(n3247), .OUT(n3251) );
  NOR2 U5237 ( .A(n3250), .B(n4400), .OUT(n6155) );
  NAND2 U5238 ( .A(n4400), .B(n3250), .OUT(n3254) );
  NAND2 U5239 ( .A(n3253), .B(n6157), .OUT(n6156) );
  NOR2 U5240 ( .A(n6157), .B(n3253), .OUT(n3257) );
  NOR2 U5241 ( .A(n3256), .B(n4404), .OUT(n6158) );
  NAND2 U5242 ( .A(n4404), .B(n3256), .OUT(n3260) );
  NAND2 U5243 ( .A(n3259), .B(n6160), .OUT(n6159) );
  NOR2 U5244 ( .A(n6160), .B(n3259), .OUT(n3263) );
  NOR2 U5245 ( .A(n3262), .B(n4408), .OUT(n6161) );
  NAND2 U5246 ( .A(n4408), .B(n3262), .OUT(n3266) );
  NAND2 U5247 ( .A(n3265), .B(n6163), .OUT(n6162) );
  NOR2 U5248 ( .A(n6163), .B(n3265), .OUT(n3269) );
  NOR2 U5249 ( .A(n3268), .B(n4412), .OUT(n6164) );
  NAND2 U5250 ( .A(n4412), .B(n3268), .OUT(n3272) );
  NAND2 U5251 ( .A(n3271), .B(n6166), .OUT(n6165) );
  NOR2 U5252 ( .A(n6166), .B(n3271), .OUT(n3275) );
  NOR2 U5253 ( .A(n3274), .B(n4416), .OUT(n6167) );
  NAND2 U5254 ( .A(n4416), .B(n3274), .OUT(n3278) );
  NAND2 U5255 ( .A(n3277), .B(n6169), .OUT(n6168) );
  NOR2 U5256 ( .A(n6169), .B(n3277), .OUT(n3281) );
  NOR2 U5257 ( .A(n3280), .B(n4420), .OUT(n6170) );
  NAND2 U5258 ( .A(n4420), .B(n3280), .OUT(n3284) );
  NAND2 U5259 ( .A(n3283), .B(n6172), .OUT(n6171) );
  NOR2 U5260 ( .A(n6172), .B(n3283), .OUT(n3287) );
  NOR2 U5261 ( .A(n3286), .B(n4424), .OUT(n6173) );
  NAND2 U5262 ( .A(n4424), .B(n3286), .OUT(n3290) );
  NAND2 U5263 ( .A(n3289), .B(n6175), .OUT(n6174) );
  NOR2 U5264 ( .A(n6175), .B(n3289), .OUT(n3293) );
  NOR2 U5265 ( .A(n3292), .B(n4428), .OUT(n6176) );
  NAND2 U5266 ( .A(n4428), .B(n3292), .OUT(n3296) );
  NAND2 U5267 ( .A(\mult_49/ab[0][30] ), .B(n6178), .OUT(n6177) );
  NOR2 U5268 ( .A(n6178), .B(\mult_49/ab[0][30] ), .OUT(n3299) );
  INV U5269 ( .IN(n3298), .OUT(n5157) );
  NAND2 U5270 ( .A(n1774), .B(n1777), .OUT(n4432) );
  NAND2 U5271 ( .A(\mult_49/ab[2][28] ), .B(n5070), .OUT(n4431) );
  NOR2 U5272 ( .A(n3298), .B(n4430), .OUT(n6179) );
  NAND2 U5273 ( .A(n4430), .B(n3298), .OUT(n3302) );
  NOR2 U5274 ( .A(n6180), .B(n4433), .OUT(n3306) );
  NOR2 U5275 ( .A(n6181), .B(n3301), .OUT(n3305) );
  NOR2 U5276 ( .A(n3304), .B(n4436), .OUT(n6182) );
  NAND2 U5277 ( .A(n4436), .B(n3304), .OUT(n3308) );
  NAND2 U5278 ( .A(n3307), .B(n6184), .OUT(n6183) );
  NOR2 U5279 ( .A(n6184), .B(n3307), .OUT(n3311) );
  NOR2 U5280 ( .A(n3310), .B(n4442), .OUT(n6185) );
  NAND2 U5281 ( .A(n4442), .B(n3310), .OUT(n3314) );
  NAND2 U5282 ( .A(n3313), .B(n6187), .OUT(n6186) );
  NOR2 U5283 ( .A(n6187), .B(n3313), .OUT(n3317) );
  NOR2 U5284 ( .A(n3316), .B(n4448), .OUT(n6188) );
  NAND2 U5285 ( .A(n4448), .B(n3316), .OUT(n3320) );
  NAND2 U5286 ( .A(n3319), .B(n6190), .OUT(n6189) );
  NOR2 U5287 ( .A(n6190), .B(n3319), .OUT(n3323) );
  NOR2 U5288 ( .A(n3322), .B(n4454), .OUT(n6191) );
  NAND2 U5289 ( .A(n4454), .B(n3322), .OUT(n3326) );
  NAND2 U5290 ( .A(n3325), .B(n6193), .OUT(n6192) );
  NOR2 U5291 ( .A(n6193), .B(n3325), .OUT(n3329) );
  NOR2 U5292 ( .A(n3328), .B(n4460), .OUT(n6194) );
  NAND2 U5293 ( .A(n4460), .B(n3328), .OUT(n3332) );
  NAND2 U5294 ( .A(n3331), .B(n6196), .OUT(n6195) );
  NOR2 U5295 ( .A(n6196), .B(n3331), .OUT(n3335) );
  NOR2 U5296 ( .A(n3334), .B(n4466), .OUT(n6197) );
  NAND2 U5297 ( .A(n4466), .B(n3334), .OUT(n3338) );
  NAND2 U5298 ( .A(n3337), .B(n6199), .OUT(n6198) );
  NOR2 U5299 ( .A(n6199), .B(n3337), .OUT(n3341) );
  NOR2 U5300 ( .A(n3340), .B(n4472), .OUT(n6200) );
  NAND2 U5301 ( .A(n4472), .B(n3340), .OUT(n3344) );
  NAND2 U5302 ( .A(n3343), .B(n6202), .OUT(n6201) );
  NOR2 U5303 ( .A(n6202), .B(n3343), .OUT(n3347) );
  NOR2 U5304 ( .A(n3346), .B(n4478), .OUT(n6203) );
  NAND2 U5305 ( .A(n4478), .B(n3346), .OUT(n3350) );
  NAND2 U5306 ( .A(n3349), .B(n6205), .OUT(n6204) );
  NOR2 U5307 ( .A(n6205), .B(n3349), .OUT(n3353) );
  NOR2 U5308 ( .A(n3352), .B(n4484), .OUT(n6206) );
  NAND2 U5309 ( .A(n4484), .B(n3352), .OUT(n3356) );
  NAND2 U5310 ( .A(n3355), .B(n6208), .OUT(n6207) );
  NOR2 U5311 ( .A(n6208), .B(n3355), .OUT(n3359) );
  NOR2 U5312 ( .A(n3358), .B(n4490), .OUT(n6209) );
  NAND2 U5313 ( .A(n4490), .B(n3358), .OUT(n3362) );
  NAND2 U5314 ( .A(n3361), .B(n6211), .OUT(n6210) );
  NOR2 U5315 ( .A(n6211), .B(n3361), .OUT(n3365) );
  NOR2 U5316 ( .A(n3364), .B(n4496), .OUT(n6212) );
  NAND2 U5317 ( .A(n4496), .B(n3364), .OUT(n3368) );
  NAND2 U5318 ( .A(n3367), .B(n6214), .OUT(n6213) );
  NOR2 U5319 ( .A(n6214), .B(n3367), .OUT(n3371) );
  NOR2 U5320 ( .A(n3370), .B(n4502), .OUT(n6215) );
  NAND2 U5321 ( .A(n4502), .B(n3370), .OUT(n3374) );
  NAND2 U5322 ( .A(n3373), .B(n6217), .OUT(n6216) );
  NOR2 U5323 ( .A(n6217), .B(n3373), .OUT(n3377) );
  NAND2 U5324 ( .A(\mult_49/ab[25][6] ), .B(n6219), .OUT(n6218) );
  NOR2 U5325 ( .A(n6219), .B(\mult_49/ab[25][6] ), .OUT(n4713) );
  INV U5326 ( .IN(n4712), .OUT(n6220) );
  NAND2 U5327 ( .A(\mult_49/ab[27][4] ), .B(n4792), .OUT(n6221) );
  NOR2 U5328 ( .A(n4792), .B(\mult_49/ab[27][4] ), .OUT(n4716) );
  NAND2 U5329 ( .A(n6220), .B(n4715), .OUT(n6222) );
  NOR2 U5330 ( .A(n4715), .B(n6220), .OUT(n4719) );
  INV U5331 ( .IN(n4718), .OUT(n6223) );
  NAND2 U5332 ( .A(\mult_49/ab[24][7] ), .B(n6225), .OUT(n6224) );
  NOR2 U5333 ( .A(n6225), .B(\mult_49/ab[24][7] ), .OUT(n4698) );
  INV U5334 ( .IN(n4697), .OUT(n6226) );
  NAND2 U5335 ( .A(n6228), .B(n4796), .OUT(n6227) );
  NOR2 U5336 ( .A(n4796), .B(n6228), .OUT(n4701) );
  NAND2 U5337 ( .A(n6226), .B(n4700), .OUT(n6229) );
  NOR2 U5338 ( .A(n4700), .B(n6226), .OUT(n4704) );
  INV U5339 ( .IN(n4703), .OUT(n6230) );
  NAND2 U5340 ( .A(\mult_49/ab[17][14] ), .B(n6232), .OUT(n6231) );
  NOR2 U5341 ( .A(n6232), .B(\mult_49/ab[17][14] ), .OUT(n4680) );
  INV U5342 ( .IN(n4679), .OUT(n6233) );
  NAND2 U5343 ( .A(\mult_49/ab[19][12] ), .B(n4798), .OUT(n6234) );
  NOR2 U5344 ( .A(n4798), .B(\mult_49/ab[19][12] ), .OUT(n4683) );
  NAND2 U5345 ( .A(n6233), .B(n4682), .OUT(n6235) );
  NOR2 U5346 ( .A(n4682), .B(n6233), .OUT(n4686) );
  INV U5347 ( .IN(n4685), .OUT(n6236) );
  NAND2 U5348 ( .A(n6238), .B(n4802), .OUT(n6237) );
  NOR2 U5349 ( .A(n4802), .B(n6238), .OUT(n4689) );
  INV U5350 ( .IN(n4688), .OUT(n6239) );
  NAND2 U5351 ( .A(\mult_49/ab[16][15] ), .B(n6241), .OUT(n6240) );
  NOR2 U5352 ( .A(n6241), .B(\mult_49/ab[16][15] ), .OUT(n4659) );
  INV U5353 ( .IN(n4658), .OUT(n6242) );
  NAND2 U5354 ( .A(n6244), .B(n4806), .OUT(n6243) );
  NOR2 U5355 ( .A(n4806), .B(n6244), .OUT(n4662) );
  NAND2 U5356 ( .A(n6242), .B(n4661), .OUT(n6245) );
  NOR2 U5357 ( .A(n4661), .B(n6242), .OUT(n4665) );
  INV U5358 ( .IN(n4664), .OUT(n6246) );
  NAND2 U5359 ( .A(\mult_49/ab[9][22] ), .B(n6248), .OUT(n6247) );
  NOR2 U5360 ( .A(n6248), .B(\mult_49/ab[9][22] ), .OUT(n4641) );
  INV U5361 ( .IN(n4640), .OUT(n6249) );
  NAND2 U5362 ( .A(\mult_49/ab[11][20] ), .B(n4808), .OUT(n6250) );
  NOR2 U5363 ( .A(n4808), .B(\mult_49/ab[11][20] ), .OUT(n4644) );
  NAND2 U5364 ( .A(n6249), .B(n4643), .OUT(n6251) );
  NOR2 U5365 ( .A(n4643), .B(n6249), .OUT(n4647) );
  INV U5366 ( .IN(n4646), .OUT(n6252) );
  NAND2 U5367 ( .A(n6254), .B(n4812), .OUT(n6253) );
  NOR2 U5368 ( .A(n4812), .B(n6254), .OUT(n4650) );
  INV U5369 ( .IN(n4649), .OUT(n6255) );
  NAND2 U5370 ( .A(\mult_49/ab[8][23] ), .B(n6257), .OUT(n6256) );
  NOR2 U5371 ( .A(n6257), .B(\mult_49/ab[8][23] ), .OUT(n4620) );
  INV U5372 ( .IN(n4619), .OUT(n6258) );
  NAND2 U5373 ( .A(n6260), .B(n4816), .OUT(n6259) );
  NOR2 U5374 ( .A(n4816), .B(n6260), .OUT(n4623) );
  NAND2 U5375 ( .A(n6258), .B(n4622), .OUT(n6261) );
  NOR2 U5376 ( .A(n4622), .B(n6258), .OUT(n4626) );
  INV U5377 ( .IN(n4625), .OUT(n6262) );
  NAND2 U5378 ( .A(\mult_49/ab[5][26] ), .B(n6264), .OUT(n6263) );
  NOR2 U5379 ( .A(n6264), .B(\mult_49/ab[5][26] ), .OUT(n4605) );
  INV U5380 ( .IN(n4604), .OUT(n6265) );
  NAND2 U5381 ( .A(\mult_49/ab[7][24] ), .B(n4818), .OUT(n6266) );
  NOR2 U5382 ( .A(n4818), .B(\mult_49/ab[7][24] ), .OUT(n4608) );
  NAND2 U5383 ( .A(n6265), .B(n4607), .OUT(n6267) );
  NOR2 U5384 ( .A(n4607), .B(n6265), .OUT(n4611) );
  INV U5385 ( .IN(n4610), .OUT(n6268) );
  NAND2 U5386 ( .A(\mult_49/ab[0][31] ), .B(n6270), .OUT(n6269) );
  NOR2 U5387 ( .A(n6270), .B(\mult_49/ab[0][31] ), .OUT(n4587) );
  INV U5388 ( .IN(n4586), .OUT(n6271) );
  NOR2 U5389 ( .A(n4820), .B(\mult_49/ab[2][29] ), .OUT(n4591) );
  NAND2 U5390 ( .A(\mult_49/ab[2][29] ), .B(n4820), .OUT(n6272) );
  NAND2 U5391 ( .A(n6271), .B(n4589), .OUT(n6273) );
  NOR2 U5392 ( .A(n4589), .B(n6271), .OUT(n4593) );
  INV U5393 ( .IN(n4592), .OUT(n6274) );
  NAND2 U5394 ( .A(\mult_49/ab[3][28] ), .B(n6276), .OUT(n6275) );
  NOR2 U5395 ( .A(n6276), .B(\mult_49/ab[3][28] ), .OUT(n4596) );
  INV U5396 ( .IN(n4595), .OUT(n6277) );
  NAND2 U5397 ( .A(n6279), .B(n4824), .OUT(n6278) );
  NOR2 U5398 ( .A(n4824), .B(n6279), .OUT(n4599) );
  NAND2 U5399 ( .A(n6277), .B(n4598), .OUT(n6280) );
  NOR2 U5400 ( .A(n4598), .B(n6277), .OUT(n4602) );
  NAND2 U5401 ( .A(n6274), .B(n4601), .OUT(n6281) );
  NOR2 U5402 ( .A(n4601), .B(n6274), .OUT(n3380) );
  INV U5403 ( .IN(n3379), .OUT(n6282) );
  NAND2 U5404 ( .A(n6284), .B(n4828), .OUT(n6283) );
  NOR2 U5405 ( .A(n4828), .B(n6284), .OUT(n4614) );
  NAND2 U5406 ( .A(n6282), .B(n4613), .OUT(n6285) );
  NOR2 U5407 ( .A(n4613), .B(n6282), .OUT(n4617) );
  NAND2 U5408 ( .A(n6268), .B(n4616), .OUT(n6286) );
  NOR2 U5409 ( .A(n4616), .B(n6268), .OUT(n3383) );
  INV U5410 ( .IN(n3382), .OUT(n6287) );
  NAND2 U5411 ( .A(n6289), .B(n4832), .OUT(n6288) );
  NOR2 U5412 ( .A(n4832), .B(n6289), .OUT(n4629) );
  NAND2 U5413 ( .A(n6287), .B(n4628), .OUT(n6290) );
  NOR2 U5414 ( .A(n4628), .B(n6287), .OUT(n4632) );
  NAND2 U5415 ( .A(n6262), .B(n4631), .OUT(n6291) );
  NOR2 U5416 ( .A(n4631), .B(n6262), .OUT(n3386) );
  INV U5417 ( .IN(n3385), .OUT(n6292) );
  NAND2 U5418 ( .A(\mult_49/ab[13][18] ), .B(n6294), .OUT(n6293) );
  NOR2 U5419 ( .A(n6294), .B(\mult_49/ab[13][18] ), .OUT(n4635) );
  INV U5420 ( .IN(n4634), .OUT(n6295) );
  NAND2 U5421 ( .A(\mult_49/ab[15][16] ), .B(n4834), .OUT(n6296) );
  NOR2 U5422 ( .A(n4834), .B(\mult_49/ab[15][16] ), .OUT(n4638) );
  NAND2 U5423 ( .A(n6295), .B(n4637), .OUT(n6297) );
  NOR2 U5424 ( .A(n4637), .B(n6295), .OUT(n3389) );
  NAND2 U5425 ( .A(n6292), .B(n3388), .OUT(n6298) );
  NOR2 U5426 ( .A(n3388), .B(n6292), .OUT(n4653) );
  NAND2 U5427 ( .A(n6255), .B(n4652), .OUT(n6299) );
  NOR2 U5428 ( .A(n4652), .B(n6255), .OUT(n4656) );
  NAND2 U5429 ( .A(n6252), .B(n4655), .OUT(n6300) );
  NOR2 U5430 ( .A(n4655), .B(n6252), .OUT(n3392) );
  INV U5431 ( .IN(n3391), .OUT(n6301) );
  NAND2 U5432 ( .A(n6303), .B(n4838), .OUT(n6302) );
  NOR2 U5433 ( .A(n4838), .B(n6303), .OUT(n4668) );
  NAND2 U5434 ( .A(n6301), .B(n4667), .OUT(n6304) );
  NOR2 U5435 ( .A(n4667), .B(n6301), .OUT(n4671) );
  NAND2 U5436 ( .A(n6246), .B(n4670), .OUT(n6305) );
  NOR2 U5437 ( .A(n4670), .B(n6246), .OUT(n3395) );
  INV U5438 ( .IN(n3394), .OUT(n6306) );
  NAND2 U5439 ( .A(\mult_49/ab[21][10] ), .B(n6308), .OUT(n6307) );
  NOR2 U5440 ( .A(n6308), .B(\mult_49/ab[21][10] ), .OUT(n4674) );
  INV U5441 ( .IN(n4673), .OUT(n6309) );
  NAND2 U5442 ( .A(\mult_49/ab[23][8] ), .B(n4840), .OUT(n6310) );
  NOR2 U5443 ( .A(n4840), .B(\mult_49/ab[23][8] ), .OUT(n4677) );
  NAND2 U5444 ( .A(n6309), .B(n4676), .OUT(n6311) );
  NOR2 U5445 ( .A(n4676), .B(n6309), .OUT(n3398) );
  NAND2 U5446 ( .A(n6306), .B(n3397), .OUT(n6312) );
  NOR2 U5447 ( .A(n3397), .B(n6306), .OUT(n4692) );
  NAND2 U5448 ( .A(n6239), .B(n4691), .OUT(n6313) );
  NOR2 U5449 ( .A(n4691), .B(n6239), .OUT(n4695) );
  NAND2 U5450 ( .A(n6236), .B(n4694), .OUT(n6314) );
  NOR2 U5451 ( .A(n4694), .B(n6236), .OUT(n3401) );
  INV U5452 ( .IN(n3400), .OUT(n6315) );
  NAND2 U5453 ( .A(n6317), .B(n4844), .OUT(n6316) );
  NOR2 U5454 ( .A(n4844), .B(n6317), .OUT(n4707) );
  NAND2 U5455 ( .A(n6315), .B(n4706), .OUT(n6318) );
  NOR2 U5456 ( .A(n4706), .B(n6315), .OUT(n4710) );
  NAND2 U5457 ( .A(n6230), .B(n4709), .OUT(n6319) );
  NOR2 U5458 ( .A(n4709), .B(n6230), .OUT(n3404) );
  INV U5459 ( .IN(n3403), .OUT(n6320) );
  NOR2 U5460 ( .A(n2377), .B(n4508), .OUT(n6321) );
  NAND2 U5461 ( .A(n4508), .B(n2377), .OUT(n3407) );
  NAND2 U5462 ( .A(n2407), .B(n6323), .OUT(n6322) );
  NOR2 U5463 ( .A(n6323), .B(n2407), .OUT(n3413) );
  NOR2 U5464 ( .A(n2440), .B(n4512), .OUT(n6324) );
  NAND2 U5465 ( .A(n4512), .B(n2440), .OUT(n3419) );
  NAND2 U5466 ( .A(n2476), .B(n6326), .OUT(n6325) );
  NOR2 U5467 ( .A(n6326), .B(n2476), .OUT(n3425) );
  NOR2 U5468 ( .A(n2515), .B(n4516), .OUT(n6327) );
  NAND2 U5469 ( .A(n4516), .B(n2515), .OUT(n3431) );
  NAND2 U5470 ( .A(n2557), .B(n6329), .OUT(n6328) );
  NOR2 U5471 ( .A(n6329), .B(n2557), .OUT(n3437) );
  NOR2 U5472 ( .A(n2602), .B(n4520), .OUT(n6330) );
  NAND2 U5473 ( .A(n4520), .B(n2602), .OUT(n3443) );
  NAND2 U5474 ( .A(n2650), .B(n6332), .OUT(n6331) );
  NOR2 U5475 ( .A(n6332), .B(n2650), .OUT(n3449) );
  NOR2 U5476 ( .A(n2701), .B(n4524), .OUT(n6333) );
  NAND2 U5477 ( .A(n4524), .B(n2701), .OUT(n3455) );
  NAND2 U5478 ( .A(n2755), .B(n6335), .OUT(n6334) );
  NOR2 U5479 ( .A(n6335), .B(n2755), .OUT(n3461) );
  NOR2 U5480 ( .A(n2812), .B(n4528), .OUT(n6336) );
  NAND2 U5481 ( .A(n4528), .B(n2812), .OUT(n3467) );
  NAND2 U5482 ( .A(n2872), .B(n6338), .OUT(n6337) );
  NOR2 U5483 ( .A(n6338), .B(n2872), .OUT(n3473) );
  NOR2 U5484 ( .A(n2935), .B(n4532), .OUT(n6339) );
  NAND2 U5485 ( .A(n4532), .B(n2935), .OUT(n3479) );
  NAND2 U5486 ( .A(n3001), .B(n6341), .OUT(n6340) );
  NOR2 U5487 ( .A(n6341), .B(n3001), .OUT(n3485) );
  NOR2 U5488 ( .A(n3070), .B(n4536), .OUT(n6342) );
  NAND2 U5489 ( .A(n4536), .B(n3070), .OUT(n3491) );
  NAND2 U5490 ( .A(n3142), .B(n6344), .OUT(n6343) );
  NOR2 U5491 ( .A(n6344), .B(n3142), .OUT(n3497) );
  NOR2 U5492 ( .A(n3217), .B(n4540), .OUT(n6345) );
  NAND2 U5493 ( .A(n4540), .B(n3217), .OUT(n3503) );
  NAND2 U5494 ( .A(n3295), .B(n6347), .OUT(n6346) );
  NOR2 U5495 ( .A(n6347), .B(n3295), .OUT(n3509) );
  NOR2 U5496 ( .A(n3376), .B(n4544), .OUT(n6348) );
  NAND2 U5497 ( .A(n4544), .B(n3376), .OUT(n3515) );
  NAND2 U5498 ( .A(n3406), .B(n6350), .OUT(n6349) );
  NOR2 U5499 ( .A(n6350), .B(n3406), .OUT(n3410) );
  NOR2 U5500 ( .A(n3412), .B(n4549), .OUT(n3417) );
  NAND2 U5501 ( .A(n4549), .B(n3412), .OUT(n6351) );
  INV U5502 ( .IN(n3415), .OUT(n5522) );
  NAND2 U5503 ( .A(n3418), .B(n6353), .OUT(n6352) );
  NOR2 U5504 ( .A(n6353), .B(n3418), .OUT(n3422) );
  NOR2 U5505 ( .A(n3424), .B(n4553), .OUT(n3429) );
  NAND2 U5506 ( .A(n4553), .B(n3424), .OUT(n6354) );
  INV U5507 ( .IN(n3427), .OUT(n5525) );
  NAND2 U5508 ( .A(n3430), .B(n6356), .OUT(n6355) );
  NOR2 U5509 ( .A(n6356), .B(n3430), .OUT(n3434) );
  NOR2 U5510 ( .A(n3436), .B(n4557), .OUT(n3441) );
  NAND2 U5511 ( .A(n4557), .B(n3436), .OUT(n6357) );
  INV U5512 ( .IN(n3439), .OUT(n5528) );
  NAND2 U5513 ( .A(n3442), .B(n6359), .OUT(n6358) );
  NOR2 U5514 ( .A(n6359), .B(n3442), .OUT(n3446) );
  NOR2 U5515 ( .A(n3448), .B(n4561), .OUT(n3453) );
  NAND2 U5516 ( .A(n4561), .B(n3448), .OUT(n6360) );
  INV U5517 ( .IN(n3451), .OUT(n5531) );
  NAND2 U5518 ( .A(n3454), .B(n6362), .OUT(n6361) );
  NOR2 U5519 ( .A(n6362), .B(n3454), .OUT(n3458) );
  NOR2 U5520 ( .A(n3460), .B(n4565), .OUT(n3465) );
  NAND2 U5521 ( .A(n4565), .B(n3460), .OUT(n6363) );
  INV U5522 ( .IN(n3463), .OUT(n5534) );
  NAND2 U5523 ( .A(n3466), .B(n6365), .OUT(n6364) );
  NOR2 U5524 ( .A(n6365), .B(n3466), .OUT(n3470) );
  NOR2 U5525 ( .A(n3472), .B(n4569), .OUT(n3477) );
  NAND2 U5526 ( .A(n4569), .B(n3472), .OUT(n6366) );
  INV U5527 ( .IN(n3475), .OUT(n5537) );
  NAND2 U5528 ( .A(n3478), .B(n6368), .OUT(n6367) );
  NOR2 U5529 ( .A(n6368), .B(n3478), .OUT(n3482) );
  NOR2 U5530 ( .A(n3484), .B(n4573), .OUT(n3489) );
  NAND2 U5531 ( .A(n4573), .B(n3484), .OUT(n6369) );
  INV U5532 ( .IN(n3487), .OUT(n5540) );
  NAND2 U5533 ( .A(n3490), .B(n6371), .OUT(n6370) );
  NOR2 U5534 ( .A(n6371), .B(n3490), .OUT(n3494) );
  NOR2 U5535 ( .A(n3496), .B(n4577), .OUT(n3501) );
  NAND2 U5536 ( .A(n4577), .B(n3496), .OUT(n6372) );
  INV U5537 ( .IN(n3499), .OUT(n5543) );
  NAND2 U5538 ( .A(n3502), .B(n6374), .OUT(n6373) );
  NOR2 U5539 ( .A(n6374), .B(n3502), .OUT(n3506) );
  NOR2 U5540 ( .A(n3508), .B(n4581), .OUT(n3513) );
  NAND2 U5541 ( .A(n4581), .B(n3508), .OUT(n6375) );
  INV U5542 ( .IN(n3511), .OUT(n5546) );
  NAND2 U5543 ( .A(n3514), .B(n6377), .OUT(n6376) );
  NOR2 U5544 ( .A(n6377), .B(n3514), .OUT(n3518) );
  NAND2 U5545 ( .A(n6379), .B(n4848), .OUT(n6378) );
  NOR2 U5546 ( .A(n4848), .B(n6379), .OUT(n4722) );
  NAND2 U5547 ( .A(n6320), .B(n4721), .OUT(n6380) );
  NOR2 U5548 ( .A(n4721), .B(n6320), .OUT(n4725) );
  NAND2 U5549 ( .A(n6223), .B(n4724), .OUT(n3522) );
  NOR2 U5550 ( .A(n4724), .B(n6223), .OUT(n6381) );
  NOR2 U5551 ( .A(n4850), .B(n3520), .OUT(n4735) );
  NAND2 U5552 ( .A(n3520), .B(n4850), .OUT(n6382) );
  NAND2 U5553 ( .A(\mult_49/ab[30][0] ), .B(n2027), .OUT(n4738) );
  NAND2 U5554 ( .A(n5547), .B(n2030), .OUT(n4737) );
  NOR2 U5555 ( .A(n3517), .B(n4736), .OUT(n6383) );
  NAND2 U5556 ( .A(n4736), .B(n3517), .OUT(n3523) );
  NAND2 U5557 ( .A(\mult_49/ab[29][0] ), .B(n2023), .OUT(n2028) );
  NAND2 U5558 ( .A(n5545), .B(n2026), .OUT(n4740) );
  NAND2 U5559 ( .A(\mult_49/ab[28][0] ), .B(n2019), .OUT(n2024) );
  NAND2 U5560 ( .A(n5544), .B(n2022), .OUT(n4742) );
  NOR2 U5561 ( .A(n3505), .B(n4741), .OUT(n6384) );
  NAND2 U5562 ( .A(n4741), .B(n3505), .OUT(n3525) );
  NAND2 U5563 ( .A(\mult_49/ab[27][0] ), .B(n2015), .OUT(n2020) );
  NAND2 U5564 ( .A(n5542), .B(n2018), .OUT(n4744) );
  NAND2 U5565 ( .A(\mult_49/ab[26][0] ), .B(n2011), .OUT(n2016) );
  NAND2 U5566 ( .A(n5541), .B(n2014), .OUT(n4746) );
  NOR2 U5567 ( .A(n3493), .B(n4745), .OUT(n6385) );
  NAND2 U5568 ( .A(n4745), .B(n3493), .OUT(n3527) );
  NAND2 U5569 ( .A(\mult_49/ab[25][0] ), .B(n2007), .OUT(n2012) );
  NAND2 U5570 ( .A(n5539), .B(n2010), .OUT(n4748) );
  NAND2 U5571 ( .A(\mult_49/ab[24][0] ), .B(n2003), .OUT(n2008) );
  NAND2 U5572 ( .A(n5538), .B(n2006), .OUT(n4750) );
  NOR2 U5573 ( .A(n3481), .B(n4749), .OUT(n6386) );
  NAND2 U5574 ( .A(n4749), .B(n3481), .OUT(n3529) );
  NAND2 U5575 ( .A(\mult_49/ab[23][0] ), .B(n1999), .OUT(n2004) );
  NAND2 U5576 ( .A(n5536), .B(n2002), .OUT(n4752) );
  NAND2 U5577 ( .A(\mult_49/ab[22][0] ), .B(n1995), .OUT(n2000) );
  NAND2 U5578 ( .A(n5535), .B(n1998), .OUT(n4754) );
  NOR2 U5579 ( .A(n3469), .B(n4753), .OUT(n6387) );
  NAND2 U5580 ( .A(n4753), .B(n3469), .OUT(n3531) );
  NAND2 U5581 ( .A(\mult_49/ab[3][0] ), .B(n475), .OUT(n480) );
  NAND2 U5582 ( .A(n5144), .B(n478), .OUT(n4756) );
  NAND2 U5583 ( .A(\mult_49/ab[21][0] ), .B(n1991), .OUT(n1996) );
  NAND2 U5584 ( .A(n5533), .B(n1994), .OUT(n4758) );
  NAND2 U5585 ( .A(\mult_49/ab[20][0] ), .B(n1987), .OUT(n1992) );
  NAND2 U5586 ( .A(n5532), .B(n1990), .OUT(n4760) );
  NOR2 U5587 ( .A(n3457), .B(n4759), .OUT(n6388) );
  NAND2 U5588 ( .A(n4759), .B(n3457), .OUT(n3533) );
  NAND2 U5589 ( .A(\mult_49/ab[19][0] ), .B(n1983), .OUT(n1988) );
  NAND2 U5590 ( .A(n5530), .B(n1986), .OUT(n4762) );
  NAND2 U5591 ( .A(\mult_49/ab[18][0] ), .B(n1979), .OUT(n1984) );
  NAND2 U5592 ( .A(n5529), .B(n1982), .OUT(n4764) );
  NOR2 U5593 ( .A(n3445), .B(n4763), .OUT(n6389) );
  NAND2 U5594 ( .A(n4763), .B(n3445), .OUT(n3535) );
  NAND2 U5595 ( .A(\mult_49/ab[17][0] ), .B(n1975), .OUT(n1980) );
  NAND2 U5596 ( .A(n5527), .B(n1978), .OUT(n4766) );
  NAND2 U5597 ( .A(\mult_49/ab[16][0] ), .B(n1971), .OUT(n1976) );
  NAND2 U5598 ( .A(n5526), .B(n1974), .OUT(n4768) );
  NOR2 U5599 ( .A(n3433), .B(n4767), .OUT(n6390) );
  NAND2 U5600 ( .A(n4767), .B(n3433), .OUT(n3537) );
  NAND2 U5601 ( .A(\mult_49/ab[15][0] ), .B(n1967), .OUT(n1972) );
  NAND2 U5602 ( .A(n5524), .B(n1970), .OUT(n4770) );
  NAND2 U5603 ( .A(\mult_49/ab[14][0] ), .B(n1963), .OUT(n1968) );
  NAND2 U5604 ( .A(n5523), .B(n1966), .OUT(n4772) );
  NOR2 U5605 ( .A(n3421), .B(n4771), .OUT(n6391) );
  NAND2 U5606 ( .A(n4771), .B(n3421), .OUT(n3539) );
  NAND2 U5607 ( .A(\mult_49/ab[13][0] ), .B(n1959), .OUT(n1964) );
  NAND2 U5608 ( .A(n5521), .B(n1962), .OUT(n4774) );
  NAND2 U5609 ( .A(\mult_49/ab[12][0] ), .B(n1955), .OUT(n1960) );
  NAND2 U5610 ( .A(n5520), .B(n1958), .OUT(n4776) );
  NOR2 U5611 ( .A(n3409), .B(n4775), .OUT(n6392) );
  NAND2 U5612 ( .A(n4775), .B(n3409), .OUT(n3541) );
  NAND2 U5613 ( .A(n472), .B(n471), .OUT(n4779) );
  NAND2 U5614 ( .A(\mult_49/ab[2][0] ), .B(n5098), .OUT(n4778) );
  NAND2 U5615 ( .A(n2318), .B(n6393), .OUT(n3544) );
  NOR2 U5616 ( .A(n6393), .B(n2318), .OUT(n6394) );
  NAND2 U5617 ( .A(A[9]), .B(n2032), .OUT(n3547) );
  NAND2 U5618 ( .A(B[9]), .B(n2031), .OUT(n3546) );
  INV U5619 ( .IN(n3545), .OUT(\gt_48/AEQB [9]) );
  NAND2 U5620 ( .A(A[8]), .B(n2034), .OUT(n3550) );
  NAND2 U5621 ( .A(B[8]), .B(n2033), .OUT(n3549) );
  INV U5622 ( .IN(n3548), .OUT(\gt_48/AEQB [8]) );
  NAND2 U5623 ( .A(A[7]), .B(n2036), .OUT(n3553) );
  NAND2 U5624 ( .A(B[7]), .B(n2035), .OUT(n3552) );
  INV U5625 ( .IN(n3551), .OUT(\gt_48/AEQB [7]) );
  NAND2 U5626 ( .A(A[6]), .B(n2038), .OUT(n3556) );
  NAND2 U5627 ( .A(B[6]), .B(n2037), .OUT(n3555) );
  INV U5628 ( .IN(n3554), .OUT(\gt_48/AEQB [6]) );
  NAND2 U5629 ( .A(A[5]), .B(n2040), .OUT(n3559) );
  NAND2 U5630 ( .A(B[5]), .B(n2039), .OUT(n3558) );
  INV U5631 ( .IN(n3557), .OUT(\gt_48/AEQB [5]) );
  NAND2 U5632 ( .A(A[4]), .B(n2042), .OUT(n3562) );
  NAND2 U5633 ( .A(B[4]), .B(n2041), .OUT(n3561) );
  INV U5634 ( .IN(n3560), .OUT(\gt_48/AEQB [4]) );
  NAND2 U5635 ( .A(A[3]), .B(n2044), .OUT(n3565) );
  NAND2 U5636 ( .A(B[3]), .B(n2043), .OUT(n3564) );
  INV U5637 ( .IN(n3563), .OUT(\gt_48/AEQB [3]) );
  NAND2 U5638 ( .A(\gt_48/SB ), .B(n6396), .OUT(n6395) );
  NOR2 U5639 ( .A(n6396), .B(\gt_48/SB ), .OUT(n3566) );
  INV U5640 ( .IN(\gt_48/AEQB [31]), .OUT(n4923) );
  NAND2 U5641 ( .A(A[30]), .B(n2046), .OUT(n3570) );
  NAND2 U5642 ( .A(B[30]), .B(n2045), .OUT(n3569) );
  INV U5643 ( .IN(n3568), .OUT(\gt_48/AEQB [30]) );
  NAND2 U5644 ( .A(A[2]), .B(n2048), .OUT(n3573) );
  NAND2 U5645 ( .A(B[2]), .B(n2047), .OUT(n3572) );
  INV U5646 ( .IN(n3571), .OUT(\gt_48/AEQB [2]) );
  NAND2 U5647 ( .A(A[29]), .B(n2050), .OUT(n3576) );
  NAND2 U5648 ( .A(B[29]), .B(n2049), .OUT(n3575) );
  INV U5649 ( .IN(n3574), .OUT(\gt_48/AEQB [29]) );
  NAND2 U5650 ( .A(A[28]), .B(n2052), .OUT(n3579) );
  NAND2 U5651 ( .A(B[28]), .B(n2051), .OUT(n3578) );
  INV U5652 ( .IN(n3577), .OUT(\gt_48/AEQB [28]) );
  NAND2 U5653 ( .A(A[27]), .B(n2054), .OUT(n3582) );
  NAND2 U5654 ( .A(B[27]), .B(n2053), .OUT(n3581) );
  INV U5655 ( .IN(n3580), .OUT(\gt_48/AEQB [27]) );
  NAND2 U5656 ( .A(A[26]), .B(n2056), .OUT(n3585) );
  NAND2 U5657 ( .A(B[26]), .B(n2055), .OUT(n3584) );
  INV U5658 ( .IN(n3583), .OUT(\gt_48/AEQB [26]) );
  NAND2 U5659 ( .A(A[25]), .B(n2058), .OUT(n3588) );
  NAND2 U5660 ( .A(B[25]), .B(n2057), .OUT(n3587) );
  INV U5661 ( .IN(n3586), .OUT(\gt_48/AEQB [25]) );
  NAND2 U5662 ( .A(A[24]), .B(n2060), .OUT(n3591) );
  NAND2 U5663 ( .A(B[24]), .B(n2059), .OUT(n3590) );
  INV U5664 ( .IN(n3589), .OUT(\gt_48/AEQB [24]) );
  NAND2 U5665 ( .A(A[23]), .B(n2062), .OUT(n3594) );
  NAND2 U5666 ( .A(B[23]), .B(n2061), .OUT(n3593) );
  INV U5667 ( .IN(n3592), .OUT(\gt_48/AEQB [23]) );
  NAND2 U5668 ( .A(A[22]), .B(n2064), .OUT(n3597) );
  NAND2 U5669 ( .A(B[22]), .B(n2063), .OUT(n3596) );
  INV U5670 ( .IN(n3595), .OUT(\gt_48/AEQB [22]) );
  NAND2 U5671 ( .A(A[21]), .B(n2066), .OUT(n3600) );
  NAND2 U5672 ( .A(B[21]), .B(n2065), .OUT(n3599) );
  INV U5673 ( .IN(n3598), .OUT(\gt_48/AEQB [21]) );
  NAND2 U5674 ( .A(A[20]), .B(n2068), .OUT(n3603) );
  NAND2 U5675 ( .A(B[20]), .B(n2067), .OUT(n3602) );
  INV U5676 ( .IN(n3601), .OUT(\gt_48/AEQB [20]) );
  NAND2 U5677 ( .A(A[1]), .B(n2070), .OUT(n3606) );
  NAND2 U5678 ( .A(B[1]), .B(n2069), .OUT(n3605) );
  INV U5679 ( .IN(n3604), .OUT(\gt_48/AEQB [1]) );
  NAND2 U5680 ( .A(A[19]), .B(n2072), .OUT(n3609) );
  NAND2 U5681 ( .A(B[19]), .B(n2071), .OUT(n3608) );
  INV U5682 ( .IN(n3607), .OUT(\gt_48/AEQB [19]) );
  NAND2 U5683 ( .A(A[18]), .B(n2074), .OUT(n3612) );
  NAND2 U5684 ( .A(B[18]), .B(n2073), .OUT(n3611) );
  INV U5685 ( .IN(n3610), .OUT(\gt_48/AEQB [18]) );
  NAND2 U5686 ( .A(A[17]), .B(n2076), .OUT(n3615) );
  NAND2 U5687 ( .A(B[17]), .B(n2075), .OUT(n3614) );
  INV U5688 ( .IN(n3613), .OUT(\gt_48/AEQB [17]) );
  NAND2 U5689 ( .A(A[16]), .B(n2078), .OUT(n3618) );
  NAND2 U5690 ( .A(B[16]), .B(n2077), .OUT(n3617) );
  INV U5691 ( .IN(n3616), .OUT(\gt_48/AEQB [16]) );
  NAND2 U5692 ( .A(A[15]), .B(n2080), .OUT(n3621) );
  NAND2 U5693 ( .A(B[15]), .B(n2079), .OUT(n3620) );
  INV U5694 ( .IN(n3619), .OUT(\gt_48/AEQB [15]) );
  NAND2 U5695 ( .A(A[14]), .B(n2082), .OUT(n3624) );
  NAND2 U5696 ( .A(B[14]), .B(n2081), .OUT(n3623) );
  INV U5697 ( .IN(n3622), .OUT(\gt_48/AEQB [14]) );
  NAND2 U5698 ( .A(A[13]), .B(n2084), .OUT(n3627) );
  NAND2 U5699 ( .A(B[13]), .B(n2083), .OUT(n3626) );
  INV U5700 ( .IN(n3625), .OUT(\gt_48/AEQB [13]) );
  NAND2 U5701 ( .A(A[12]), .B(n2086), .OUT(n3630) );
  NAND2 U5702 ( .A(B[12]), .B(n2085), .OUT(n3629) );
  INV U5703 ( .IN(n3628), .OUT(\gt_48/AEQB [12]) );
  NAND2 U5704 ( .A(A[11]), .B(n2088), .OUT(n3633) );
  NAND2 U5705 ( .A(B[11]), .B(n2087), .OUT(n3632) );
  INV U5706 ( .IN(n3631), .OUT(\gt_48/AEQB [11]) );
  NAND2 U5707 ( .A(A[10]), .B(n2090), .OUT(n3636) );
  NAND2 U5708 ( .A(B[10]), .B(n2089), .OUT(n3635) );
  INV U5709 ( .IN(n3634), .OUT(\gt_48/AEQB [10]) );
  NAND2 U5710 ( .A(\gt_48/AEQB [1]), .B(n2091), .OUT(n3638) );
  NAND2 U5711 ( .A(n3604), .B(n6397), .OUT(n3637) );
  NAND2 U5712 ( .A(\mult_49/ab[0][1] ), .B(n474), .OUT(n3640) );
  NAND2 U5713 ( .A(\mult_49/ab[1][0] ), .B(n473), .OUT(n3639) );
  NOR2 U5714 ( .A(n4916), .B(n4923), .OUT(n6398) );
  NAND2 U5715 ( .A(n4923), .B(n4916), .OUT(n3641) );
  NAND2 U5716 ( .A(\gt_48/AEQB [30]), .B(n5610), .OUT(n3644) );
  NAND2 U5717 ( .A(n3568), .B(n2177), .OUT(n3643) );
  NAND2 U5718 ( .A(\gt_48/AEQB [29]), .B(n5608), .OUT(n3646) );
  NAND2 U5719 ( .A(n3574), .B(n2174), .OUT(n3645) );
  NAND2 U5720 ( .A(\gt_48/AEQB [28]), .B(n5606), .OUT(n3648) );
  NAND2 U5721 ( .A(n3577), .B(n2171), .OUT(n3647) );
  NAND2 U5722 ( .A(\gt_48/AEQB [27]), .B(n5604), .OUT(n3650) );
  NAND2 U5723 ( .A(n3580), .B(n2168), .OUT(n3649) );
  NAND2 U5724 ( .A(\gt_48/AEQB [26]), .B(n5602), .OUT(n3652) );
  NAND2 U5725 ( .A(n3583), .B(n2165), .OUT(n3651) );
  NAND2 U5726 ( .A(\gt_48/AEQB [25]), .B(n5600), .OUT(n3654) );
  NAND2 U5727 ( .A(n3586), .B(n2162), .OUT(n3653) );
  NAND2 U5728 ( .A(\gt_48/AEQB [24]), .B(n5598), .OUT(n3656) );
  NAND2 U5729 ( .A(n3589), .B(n2159), .OUT(n3655) );
  NAND2 U5730 ( .A(\gt_48/AEQB [23]), .B(n5596), .OUT(n3658) );
  NAND2 U5731 ( .A(n3592), .B(n2156), .OUT(n3657) );
  NAND2 U5732 ( .A(\gt_48/AEQB [22]), .B(n5594), .OUT(n3660) );
  NAND2 U5733 ( .A(n3595), .B(n2153), .OUT(n3659) );
  NAND2 U5734 ( .A(\gt_48/AEQB [21]), .B(n5592), .OUT(n3662) );
  NAND2 U5735 ( .A(n3598), .B(n2150), .OUT(n3661) );
  NAND2 U5736 ( .A(\gt_48/AEQB [20]), .B(n5590), .OUT(n3664) );
  NAND2 U5737 ( .A(n3601), .B(n2147), .OUT(n3663) );
  NAND2 U5738 ( .A(\gt_48/AEQB [19]), .B(n5588), .OUT(n3666) );
  NAND2 U5739 ( .A(n3607), .B(n2144), .OUT(n3665) );
  NAND2 U5740 ( .A(\gt_48/AEQB [18]), .B(n5586), .OUT(n3668) );
  NAND2 U5741 ( .A(n3610), .B(n2141), .OUT(n3667) );
  NAND2 U5742 ( .A(\gt_48/AEQB [17]), .B(n5584), .OUT(n3670) );
  NAND2 U5743 ( .A(n3613), .B(n2138), .OUT(n3669) );
  NAND2 U5744 ( .A(\gt_48/AEQB [16]), .B(n5582), .OUT(n3672) );
  NAND2 U5745 ( .A(n3616), .B(n2135), .OUT(n3671) );
  NAND2 U5746 ( .A(\gt_48/AEQB [15]), .B(n5580), .OUT(n3674) );
  NAND2 U5747 ( .A(n3619), .B(n2132), .OUT(n3673) );
  NAND2 U5748 ( .A(\gt_48/AEQB [14]), .B(n5578), .OUT(n3676) );
  NAND2 U5749 ( .A(n3622), .B(n2129), .OUT(n3675) );
  NAND2 U5750 ( .A(\gt_48/AEQB [13]), .B(n5576), .OUT(n3678) );
  NAND2 U5751 ( .A(n3625), .B(n2126), .OUT(n3677) );
  NAND2 U5752 ( .A(\gt_48/AEQB [12]), .B(n5574), .OUT(n3680) );
  NAND2 U5753 ( .A(n3628), .B(n2123), .OUT(n3679) );
  NAND2 U5754 ( .A(\gt_48/AEQB [11]), .B(n5572), .OUT(n3682) );
  NAND2 U5755 ( .A(n3631), .B(n2120), .OUT(n3681) );
  NAND2 U5756 ( .A(\gt_48/AEQB [10]), .B(n5570), .OUT(n3684) );
  NAND2 U5757 ( .A(n3634), .B(n2117), .OUT(n3683) );
  NAND2 U5758 ( .A(\gt_48/AEQB [9]), .B(n5568), .OUT(n3686) );
  NAND2 U5759 ( .A(n3545), .B(n2114), .OUT(n3685) );
  NAND2 U5760 ( .A(\gt_48/AEQB [8]), .B(n5566), .OUT(n3688) );
  NAND2 U5761 ( .A(n3548), .B(n2111), .OUT(n3687) );
  NAND2 U5762 ( .A(\gt_48/AEQB [7]), .B(n5564), .OUT(n3690) );
  NAND2 U5763 ( .A(n3551), .B(n2108), .OUT(n3689) );
  NAND2 U5764 ( .A(\gt_48/AEQB [6]), .B(n5562), .OUT(n3692) );
  NAND2 U5765 ( .A(n3554), .B(n2105), .OUT(n3691) );
  NAND2 U5766 ( .A(\gt_48/AEQB [5]), .B(n5560), .OUT(n3694) );
  NAND2 U5767 ( .A(n3557), .B(n2102), .OUT(n3693) );
  NAND2 U5768 ( .A(\gt_48/AEQB [4]), .B(n5558), .OUT(n3696) );
  NAND2 U5769 ( .A(n3560), .B(n2099), .OUT(n3695) );
  NAND2 U5770 ( .A(\gt_48/AEQB [3]), .B(n5556), .OUT(n3698) );
  NAND2 U5771 ( .A(n3563), .B(n2096), .OUT(n3697) );
  NAND2 U5772 ( .A(\gt_48/AEQB [2]), .B(n5554), .OUT(n3700) );
  NAND2 U5773 ( .A(n3571), .B(n2093), .OUT(n3699) );
  NAND2 U5774 ( .A(\gt_48/AEQB [1]), .B(n2092), .OUT(n3702) );
  NAND2 U5775 ( .A(n3604), .B(n289), .OUT(n3701) );
  INV U5776 ( .IN(n5711), .OUT(n2346) );
  INV U5777 ( .IN(n5712), .OUT(n2348) );
  INV U5778 ( .IN(n5713), .OUT(n2350) );
  INV U5779 ( .IN(n5714), .OUT(n2352) );
  INV U5780 ( .IN(n4852), .OUT(n4854) );
  INV U5781 ( .IN(n6383), .OUT(n3524) );
  INV U5782 ( .IN(n6384), .OUT(n3526) );
  INV U5783 ( .IN(n6385), .OUT(n3528) );
  INV U5784 ( .IN(n6386), .OUT(n3530) );
  INV U5785 ( .IN(n6387), .OUT(n3532) );
  INV U5786 ( .IN(n6388), .OUT(n3534) );
  INV U5787 ( .IN(n6389), .OUT(n3536) );
  INV U5788 ( .IN(n6390), .OUT(n3538) );
  INV U5789 ( .IN(n6391), .OUT(n3540) );
  INV U5790 ( .IN(n6392), .OUT(n3542) );
  INV U5791 ( .IN(\mult_49/ab[0][2] ), .OUT(n437) );
  INV U5792 ( .IN(\mult_49/ab[0][3] ), .OUT(n405) );
  INV U5793 ( .IN(\mult_49/ab[0][4] ), .OUT(n377) );
  INV U5794 ( .IN(\mult_49/ab[0][5] ), .OUT(n353) );
  INV U5795 ( .IN(\mult_49/ab[0][6] ), .OUT(n333) );
  INV U5796 ( .IN(\mult_49/ab[0][7] ), .OUT(n317) );
  INV U5797 ( .IN(\mult_49/ab[0][8] ), .OUT(n305) );
  INV U5798 ( .IN(\mult_49/ab[0][9] ), .OUT(n297) );
  INV U5799 ( .IN(\mult_49/ab[0][10] ), .OUT(n292) );
  INV U5800 ( .IN(\mult_49/ab[0][11] ), .OUT(n516) );
  INV U5801 ( .IN(\mult_49/ab[0][12] ), .OUT(n552) );
  INV U5802 ( .IN(\mult_49/ab[0][13] ), .OUT(n592) );
  INV U5803 ( .IN(\mult_49/ab[0][14] ), .OUT(n636) );
  INV U5804 ( .IN(\mult_49/ab[0][15] ), .OUT(n684) );
  INV U5805 ( .IN(\mult_49/ab[0][16] ), .OUT(n736) );
  INV U5806 ( .IN(\mult_49/ab[0][17] ), .OUT(n792) );
  INV U5807 ( .IN(\mult_49/ab[0][18] ), .OUT(n852) );
  INV U5808 ( .IN(\mult_49/ab[0][19] ), .OUT(n916) );
  INV U5809 ( .IN(\mult_49/ab[0][20] ), .OUT(n984) );
  INV U5810 ( .IN(\mult_49/ab[0][21] ), .OUT(n1056) );
  INV U5811 ( .IN(\mult_49/ab[0][22] ), .OUT(n1132) );
  INV U5812 ( .IN(\mult_49/ab[0][23] ), .OUT(n1212) );
  INV U5813 ( .IN(\mult_49/ab[0][24] ), .OUT(n1296) );
  INV U5814 ( .IN(\mult_49/ab[0][25] ), .OUT(n1384) );
  INV U5815 ( .IN(\mult_49/ab[0][26] ), .OUT(n1476) );
  INV U5816 ( .IN(\mult_49/ab[0][27] ), .OUT(n1572) );
  INV U5817 ( .IN(\mult_49/ab[0][28] ), .OUT(n1672) );
  INV U5818 ( .IN(\mult_49/ab[0][29] ), .OUT(n1776) );
  INV U5819 ( .IN(n5717), .OUT(n4731) );
  INV U5820 ( .IN(n6382), .OUT(n4734) );
  INV U5821 ( .IN(\mult_49/ab[0][1] ), .OUT(n473) );
  INV U5822 ( .IN(n3703), .OUT(n5699) );
  INV U5823 ( .IN(n3706), .OUT(n5686) );
  INV U5824 ( .IN(n3709), .OUT(n5701) );
  INV U5825 ( .IN(n3711), .OUT(n5674) );
  INV U5826 ( .IN(n3714), .OUT(n5689) );
  INV U5827 ( .IN(n3718), .OUT(n5665) );
  INV U5828 ( .IN(n3721), .OUT(n5677) );
  INV U5829 ( .IN(n3727), .OUT(n5656) );
  INV U5830 ( .IN(n3730), .OUT(n5668) );
  INV U5831 ( .IN(n3738), .OUT(n5650) );
  INV U5832 ( .IN(n3741), .OUT(n5659) );
  INV U5833 ( .IN(n3751), .OUT(n5644) );
  INV U5834 ( .IN(n3754), .OUT(n5653) );
  INV U5835 ( .IN(n3766), .OUT(n5641) );
  INV U5836 ( .IN(n3769), .OUT(n5647) );
  INV U5837 ( .IN(n3783), .OUT(n5637) );
  INV U5838 ( .IN(n3786), .OUT(n5640) );
  INV U5839 ( .IN(n3818), .OUT(n5718) );
  INV U5840 ( .IN(n3821), .OUT(n5721) );
  INV U5841 ( .IN(n3835), .OUT(n5731) );
  INV U5842 ( .IN(n3838), .OUT(n5734) );
  INV U5843 ( .IN(n3854), .OUT(n5745) );
  INV U5844 ( .IN(n3857), .OUT(n5748) );
  INV U5845 ( .IN(n3875), .OUT(n5761) );
  INV U5846 ( .IN(n3878), .OUT(n5764) );
  INV U5847 ( .IN(n3898), .OUT(n5778) );
  INV U5848 ( .IN(n3901), .OUT(n5781) );
  INV U5849 ( .IN(n3923), .OUT(n5797) );
  INV U5850 ( .IN(n3926), .OUT(n5800) );
  INV U5851 ( .IN(n3950), .OUT(n5817) );
  INV U5852 ( .IN(n3953), .OUT(n5820) );
  INV U5853 ( .IN(n3979), .OUT(n5839) );
  INV U5854 ( .IN(n3982), .OUT(n5842) );
  INV U5855 ( .IN(n4010), .OUT(n5862) );
  INV U5856 ( .IN(n4013), .OUT(n5865) );
  INV U5857 ( .IN(n4043), .OUT(n5887) );
  INV U5858 ( .IN(n4046), .OUT(n5890) );
  INV U5859 ( .IN(n4078), .OUT(n5913) );
  INV U5860 ( .IN(n4081), .OUT(n5916) );
  INV U5861 ( .IN(n4115), .OUT(n5941) );
  INV U5862 ( .IN(n4118), .OUT(n5944) );
  INV U5863 ( .IN(n4154), .OUT(n5970) );
  INV U5864 ( .IN(n4157), .OUT(n5973) );
  INV U5865 ( .IN(n4195), .OUT(n6001) );
  INV U5866 ( .IN(n4198), .OUT(n6004) );
  INV U5867 ( .IN(n4238), .OUT(n6033) );
  INV U5868 ( .IN(n4241), .OUT(n6036) );
  INV U5869 ( .IN(n4283), .OUT(n6067) );
  INV U5870 ( .IN(n4286), .OUT(n6070) );
  INV U5871 ( .IN(n4330), .OUT(n6102) );
  INV U5872 ( .IN(n4333), .OUT(n6105) );
  INV U5873 ( .IN(n4379), .OUT(n6139) );
  INV U5874 ( .IN(n4382), .OUT(n6142) );
  INV U5875 ( .IN(\mult_49/ab[1][29] ), .OUT(n6178) );
  INV U5876 ( .IN(n4433), .OUT(n6181) );
  INV U5877 ( .IN(n4846), .OUT(n6379) );
  INV U5878 ( .IN(n4842), .OUT(n6317) );
  INV U5879 ( .IN(\mult_49/ab[22][9] ), .OUT(n6308) );
  INV U5880 ( .IN(n4836), .OUT(n6303) );
  INV U5881 ( .IN(\mult_49/ab[14][17] ), .OUT(n6294) );
  INV U5882 ( .IN(n4830), .OUT(n6289) );
  INV U5883 ( .IN(n4826), .OUT(n6284) );
  INV U5884 ( .IN(n4821), .OUT(n6279) );
  INV U5885 ( .IN(\mult_49/ab[4][27] ), .OUT(n6276) );
  INV U5886 ( .IN(\mult_49/ab[1][30] ), .OUT(n6270) );
  INV U5887 ( .IN(\mult_49/ab[6][25] ), .OUT(n6264) );
  INV U5888 ( .IN(n4814), .OUT(n6260) );
  INV U5889 ( .IN(\mult_49/ab[12][19] ), .OUT(n6257) );
  INV U5890 ( .IN(n4810), .OUT(n6254) );
  INV U5891 ( .IN(\mult_49/ab[10][21] ), .OUT(n6248) );
  INV U5892 ( .IN(n4804), .OUT(n6244) );
  INV U5893 ( .IN(\mult_49/ab[20][11] ), .OUT(n6241) );
  INV U5894 ( .IN(n4800), .OUT(n6238) );
  INV U5895 ( .IN(\mult_49/ab[18][13] ), .OUT(n6232) );
  INV U5896 ( .IN(n4794), .OUT(n6228) );
  INV U5897 ( .IN(\mult_49/ab[28][3] ), .OUT(n6225) );
  INV U5898 ( .IN(\mult_49/ab[26][5] ), .OUT(n6219) );
  INV U5899 ( .IN(\mult_49/ab[30][1] ), .OUT(n5716) );
  INV U5900 ( .IN(n2321), .OUT(n4869) );
  INV U5901 ( .IN(n4777), .OUT(n6393) );
  INV U5902 ( .IN(\gt_48/SA ), .OUT(n6396) );
  INV U5903 ( .IN(\mult_49/ab[1][0] ), .OUT(n474) );
  INV U5904 ( .IN(\mult_49/ab[1][1] ), .OUT(n438) );
  INV U5905 ( .IN(\mult_49/ab[1][2] ), .OUT(n406) );
  INV U5906 ( .IN(n5698), .OUT(n2323) );
  INV U5907 ( .IN(\mult_49/ab[1][3] ), .OUT(n378) );
  INV U5908 ( .IN(n5687), .OUT(n2295) );
  INV U5909 ( .IN(n2294), .OUT(n5700) );
  INV U5910 ( .IN(\mult_49/ab[1][4] ), .OUT(n354) );
  INV U5911 ( .IN(n5675), .OUT(n2271) );
  INV U5912 ( .IN(n2270), .OUT(n5688) );
  INV U5913 ( .IN(n5702), .OUT(n2328) );
  INV U5914 ( .IN(\mult_49/ab[1][5] ), .OUT(n334) );
  INV U5915 ( .IN(n5666), .OUT(n2250) );
  INV U5916 ( .IN(n2249), .OUT(n5676) );
  INV U5917 ( .IN(n5690), .OUT(n2302) );
  INV U5918 ( .IN(n3725), .OUT(n5704) );
  INV U5919 ( .IN(n5703), .OUT(n2332) );
  INV U5920 ( .IN(\mult_49/ab[1][6] ), .OUT(n318) );
  INV U5921 ( .IN(n5657), .OUT(n2232) );
  INV U5922 ( .IN(n2231), .OUT(n5667) );
  INV U5923 ( .IN(n5678), .OUT(n2278) );
  INV U5924 ( .IN(n3734), .OUT(n5692) );
  INV U5925 ( .IN(n5691), .OUT(n2305) );
  INV U5926 ( .IN(n5705), .OUT(n2334) );
  INV U5927 ( .IN(\mult_49/ab[1][7] ), .OUT(n306) );
  INV U5928 ( .IN(n5651), .OUT(n2217) );
  INV U5929 ( .IN(n2216), .OUT(n5658) );
  INV U5930 ( .IN(n5669), .OUT(n2257) );
  INV U5931 ( .IN(n3745), .OUT(n5680) );
  INV U5932 ( .IN(n5679), .OUT(n2281) );
  INV U5933 ( .IN(n5693), .OUT(n2308) );
  INV U5934 ( .IN(n3749), .OUT(n5707) );
  INV U5935 ( .IN(n5706), .OUT(n2338) );
  INV U5936 ( .IN(\mult_49/ab[1][8] ), .OUT(n298) );
  INV U5937 ( .IN(n5645), .OUT(n2205) );
  INV U5938 ( .IN(n2204), .OUT(n5652) );
  INV U5939 ( .IN(n5660), .OUT(n2239) );
  INV U5940 ( .IN(n3758), .OUT(n5671) );
  INV U5941 ( .IN(n5670), .OUT(n2260) );
  INV U5942 ( .IN(n5681), .OUT(n2284) );
  INV U5943 ( .IN(n3762), .OUT(n5695) );
  INV U5944 ( .IN(n5694), .OUT(n2311) );
  INV U5945 ( .IN(n5708), .OUT(n2340) );
  INV U5946 ( .IN(\mult_49/ab[1][9] ), .OUT(n293) );
  INV U5947 ( .IN(n5642), .OUT(n2196) );
  INV U5948 ( .IN(n2195), .OUT(n5646) );
  INV U5949 ( .IN(n5654), .OUT(n2224) );
  INV U5950 ( .IN(n3773), .OUT(n5662) );
  INV U5951 ( .IN(n5661), .OUT(n2242) );
  INV U5952 ( .IN(n5672), .OUT(n2263) );
  INV U5953 ( .IN(n3777), .OUT(n5683) );
  INV U5954 ( .IN(n5682), .OUT(n2287) );
  INV U5955 ( .IN(n5696), .OUT(n2314) );
  INV U5956 ( .IN(n3781), .OUT(n5710) );
  INV U5957 ( .IN(n5709), .OUT(n2344) );
  INV U5958 ( .IN(\mult_49/ab[1][10] ), .OUT(n515) );
  INV U5959 ( .IN(n5638), .OUT(n2184) );
  INV U5960 ( .IN(n2183), .OUT(n5639) );
  INV U5961 ( .IN(n5643), .OUT(n2200) );
  INV U5962 ( .IN(n3790), .OUT(n5649) );
  INV U5963 ( .IN(n5648), .OUT(n2212) );
  INV U5964 ( .IN(n5655), .OUT(n2227) );
  INV U5965 ( .IN(n3794), .OUT(n5664) );
  INV U5966 ( .IN(n5663), .OUT(n2245) );
  INV U5967 ( .IN(n5673), .OUT(n2266) );
  INV U5968 ( .IN(n3798), .OUT(n5685) );
  INV U5969 ( .IN(n5684), .OUT(n2290) );
  INV U5970 ( .IN(n5697), .OUT(n2316) );
  INV U5971 ( .IN(n4781), .OUT(n4782) );
  INV U5972 ( .IN(n4784), .OUT(n4785) );
  INV U5973 ( .IN(n4787), .OUT(n4788) );
  INV U5974 ( .IN(n4790), .OUT(n4791) );
  INV U5975 ( .IN(\mult_49/ab[1][11] ), .OUT(n551) );
  INV U5976 ( .IN(n5719), .OUT(n2357) );
  INV U5977 ( .IN(n2356), .OUT(n5720) );
  INV U5978 ( .IN(n5722), .OUT(n2364) );
  INV U5979 ( .IN(n3825), .OUT(n5724) );
  INV U5980 ( .IN(n5723), .OUT(n2367) );
  INV U5981 ( .IN(n5725), .OUT(n2370) );
  INV U5982 ( .IN(n3829), .OUT(n5727) );
  INV U5983 ( .IN(n5726), .OUT(n2373) );
  INV U5984 ( .IN(n5728), .OUT(n2376) );
  INV U5985 ( .IN(n3833), .OUT(n5730) );
  INV U5986 ( .IN(n5729), .OUT(n2379) );
  INV U5987 ( .IN(n6321), .OUT(n3408) );
  INV U5988 ( .IN(n4547), .OUT(n6350) );
  INV U5989 ( .IN(n6349), .OUT(n3411) );
  INV U5990 ( .IN(\mult_49/ab[1][12] ), .OUT(n591) );
  INV U5991 ( .IN(n5732), .OUT(n2384) );
  INV U5992 ( .IN(n2383), .OUT(n5733) );
  INV U5993 ( .IN(n5735), .OUT(n2391) );
  INV U5994 ( .IN(n3842), .OUT(n5737) );
  INV U5995 ( .IN(n5736), .OUT(n2394) );
  INV U5996 ( .IN(n5738), .OUT(n2397) );
  INV U5997 ( .IN(n3846), .OUT(n5740) );
  INV U5998 ( .IN(n5739), .OUT(n2400) );
  INV U5999 ( .IN(n5741), .OUT(n2403) );
  INV U6000 ( .IN(n3850), .OUT(n5743) );
  INV U6001 ( .IN(n5742), .OUT(n2406) );
  INV U6002 ( .IN(n5744), .OUT(n2409) );
  INV U6003 ( .IN(n4510), .OUT(n6323) );
  INV U6004 ( .IN(n6322), .OUT(n3414) );
  INV U6005 ( .IN(n6351), .OUT(n3416) );
  INV U6006 ( .IN(\mult_49/ab[1][13] ), .OUT(n635) );
  INV U6007 ( .IN(n5746), .OUT(n2414) );
  INV U6008 ( .IN(n2413), .OUT(n5747) );
  INV U6009 ( .IN(n5749), .OUT(n2421) );
  INV U6010 ( .IN(n3861), .OUT(n5751) );
  INV U6011 ( .IN(n5750), .OUT(n2424) );
  INV U6012 ( .IN(n5752), .OUT(n2427) );
  INV U6013 ( .IN(n3865), .OUT(n5754) );
  INV U6014 ( .IN(n5753), .OUT(n2430) );
  INV U6015 ( .IN(n5755), .OUT(n2433) );
  INV U6016 ( .IN(n3869), .OUT(n5757) );
  INV U6017 ( .IN(n5756), .OUT(n2436) );
  INV U6018 ( .IN(n5758), .OUT(n2439) );
  INV U6019 ( .IN(n3873), .OUT(n5760) );
  INV U6020 ( .IN(n5759), .OUT(n2442) );
  INV U6021 ( .IN(n6324), .OUT(n3420) );
  INV U6022 ( .IN(n4551), .OUT(n6353) );
  INV U6023 ( .IN(n6352), .OUT(n3423) );
  INV U6024 ( .IN(\mult_49/ab[1][14] ), .OUT(n683) );
  INV U6025 ( .IN(n5762), .OUT(n2447) );
  INV U6026 ( .IN(n2446), .OUT(n5763) );
  INV U6027 ( .IN(n5765), .OUT(n2454) );
  INV U6028 ( .IN(n3882), .OUT(n5767) );
  INV U6029 ( .IN(n5766), .OUT(n2457) );
  INV U6030 ( .IN(n5768), .OUT(n2460) );
  INV U6031 ( .IN(n3886), .OUT(n5770) );
  INV U6032 ( .IN(n5769), .OUT(n2463) );
  INV U6033 ( .IN(n5771), .OUT(n2466) );
  INV U6034 ( .IN(n3890), .OUT(n5773) );
  INV U6035 ( .IN(n5772), .OUT(n2469) );
  INV U6036 ( .IN(n5774), .OUT(n2472) );
  INV U6037 ( .IN(n3894), .OUT(n5776) );
  INV U6038 ( .IN(n5775), .OUT(n2475) );
  INV U6039 ( .IN(n5777), .OUT(n2478) );
  INV U6040 ( .IN(n4514), .OUT(n6326) );
  INV U6041 ( .IN(n6325), .OUT(n3426) );
  INV U6042 ( .IN(n6354), .OUT(n3428) );
  INV U6043 ( .IN(\mult_49/ab[1][15] ), .OUT(n735) );
  INV U6044 ( .IN(n5779), .OUT(n2483) );
  INV U6045 ( .IN(n2482), .OUT(n5780) );
  INV U6046 ( .IN(n5782), .OUT(n2490) );
  INV U6047 ( .IN(n3905), .OUT(n5784) );
  INV U6048 ( .IN(n5783), .OUT(n2493) );
  INV U6049 ( .IN(n5785), .OUT(n2496) );
  INV U6050 ( .IN(n3909), .OUT(n5787) );
  INV U6051 ( .IN(n5786), .OUT(n2499) );
  INV U6052 ( .IN(n5788), .OUT(n2502) );
  INV U6053 ( .IN(n3913), .OUT(n5790) );
  INV U6054 ( .IN(n5789), .OUT(n2505) );
  INV U6055 ( .IN(n5791), .OUT(n2508) );
  INV U6056 ( .IN(n3917), .OUT(n5793) );
  INV U6057 ( .IN(n5792), .OUT(n2511) );
  INV U6058 ( .IN(n5794), .OUT(n2514) );
  INV U6059 ( .IN(n3921), .OUT(n5796) );
  INV U6060 ( .IN(n5795), .OUT(n2517) );
  INV U6061 ( .IN(n6327), .OUT(n3432) );
  INV U6062 ( .IN(n4555), .OUT(n6356) );
  INV U6063 ( .IN(n6355), .OUT(n3435) );
  INV U6064 ( .IN(\mult_49/ab[1][16] ), .OUT(n791) );
  INV U6065 ( .IN(n5798), .OUT(n2522) );
  INV U6066 ( .IN(n2521), .OUT(n5799) );
  INV U6067 ( .IN(n5801), .OUT(n2529) );
  INV U6068 ( .IN(n3930), .OUT(n5803) );
  INV U6069 ( .IN(n5802), .OUT(n2532) );
  INV U6070 ( .IN(n5804), .OUT(n2535) );
  INV U6071 ( .IN(n3934), .OUT(n5806) );
  INV U6072 ( .IN(n5805), .OUT(n2538) );
  INV U6073 ( .IN(n5807), .OUT(n2541) );
  INV U6074 ( .IN(n3938), .OUT(n5809) );
  INV U6075 ( .IN(n5808), .OUT(n2544) );
  INV U6076 ( .IN(n5810), .OUT(n2547) );
  INV U6077 ( .IN(n3942), .OUT(n5812) );
  INV U6078 ( .IN(n5811), .OUT(n2550) );
  INV U6079 ( .IN(n5813), .OUT(n2553) );
  INV U6080 ( .IN(n3946), .OUT(n5815) );
  INV U6081 ( .IN(n5814), .OUT(n2556) );
  INV U6082 ( .IN(n5816), .OUT(n2559) );
  INV U6083 ( .IN(n4518), .OUT(n6329) );
  INV U6084 ( .IN(n6328), .OUT(n3438) );
  INV U6085 ( .IN(n6357), .OUT(n3440) );
  INV U6086 ( .IN(\mult_49/ab[1][17] ), .OUT(n851) );
  INV U6087 ( .IN(n5818), .OUT(n2564) );
  INV U6088 ( .IN(n2563), .OUT(n5819) );
  INV U6089 ( .IN(n5821), .OUT(n2571) );
  INV U6090 ( .IN(n3957), .OUT(n5823) );
  INV U6091 ( .IN(n5822), .OUT(n2574) );
  INV U6092 ( .IN(n5824), .OUT(n2577) );
  INV U6093 ( .IN(n3961), .OUT(n5826) );
  INV U6094 ( .IN(n5825), .OUT(n2580) );
  INV U6095 ( .IN(n5827), .OUT(n2583) );
  INV U6096 ( .IN(n3965), .OUT(n5829) );
  INV U6097 ( .IN(n5828), .OUT(n2586) );
  INV U6098 ( .IN(n5830), .OUT(n2589) );
  INV U6099 ( .IN(n3969), .OUT(n5832) );
  INV U6100 ( .IN(n5831), .OUT(n2592) );
  INV U6101 ( .IN(n5833), .OUT(n2595) );
  INV U6102 ( .IN(n3973), .OUT(n5835) );
  INV U6103 ( .IN(n5834), .OUT(n2598) );
  INV U6104 ( .IN(n5836), .OUT(n2601) );
  INV U6105 ( .IN(n3977), .OUT(n5838) );
  INV U6106 ( .IN(n5837), .OUT(n2604) );
  INV U6107 ( .IN(n6330), .OUT(n3444) );
  INV U6108 ( .IN(n4559), .OUT(n6359) );
  INV U6109 ( .IN(n6358), .OUT(n3447) );
  INV U6110 ( .IN(\mult_49/ab[1][18] ), .OUT(n915) );
  INV U6111 ( .IN(n5840), .OUT(n2609) );
  INV U6112 ( .IN(n2608), .OUT(n5841) );
  INV U6113 ( .IN(n5843), .OUT(n2616) );
  INV U6114 ( .IN(n3986), .OUT(n5845) );
  INV U6115 ( .IN(n5844), .OUT(n2619) );
  INV U6116 ( .IN(n5846), .OUT(n2622) );
  INV U6117 ( .IN(n3990), .OUT(n5848) );
  INV U6118 ( .IN(n5847), .OUT(n2625) );
  INV U6119 ( .IN(n5849), .OUT(n2628) );
  INV U6120 ( .IN(n3994), .OUT(n5851) );
  INV U6121 ( .IN(n5850), .OUT(n2631) );
  INV U6122 ( .IN(n5852), .OUT(n2634) );
  INV U6123 ( .IN(n3998), .OUT(n5854) );
  INV U6124 ( .IN(n5853), .OUT(n2637) );
  INV U6125 ( .IN(n5855), .OUT(n2640) );
  INV U6126 ( .IN(n4002), .OUT(n5857) );
  INV U6127 ( .IN(n5856), .OUT(n2643) );
  INV U6128 ( .IN(n5858), .OUT(n2646) );
  INV U6129 ( .IN(n4006), .OUT(n5860) );
  INV U6130 ( .IN(n5859), .OUT(n2649) );
  INV U6131 ( .IN(n5861), .OUT(n2652) );
  INV U6132 ( .IN(n4522), .OUT(n6332) );
  INV U6133 ( .IN(n6331), .OUT(n3450) );
  INV U6134 ( .IN(n6360), .OUT(n3452) );
  INV U6135 ( .IN(\mult_49/ab[1][19] ), .OUT(n983) );
  INV U6136 ( .IN(n5863), .OUT(n2657) );
  INV U6137 ( .IN(n2656), .OUT(n5864) );
  INV U6138 ( .IN(n5866), .OUT(n2664) );
  INV U6139 ( .IN(n4017), .OUT(n5868) );
  INV U6140 ( .IN(n5867), .OUT(n2667) );
  INV U6141 ( .IN(n5869), .OUT(n2670) );
  INV U6142 ( .IN(n4021), .OUT(n5871) );
  INV U6143 ( .IN(n5870), .OUT(n2673) );
  INV U6144 ( .IN(n5872), .OUT(n2676) );
  INV U6145 ( .IN(n4025), .OUT(n5874) );
  INV U6146 ( .IN(n5873), .OUT(n2679) );
  INV U6147 ( .IN(n5875), .OUT(n2682) );
  INV U6148 ( .IN(n4029), .OUT(n5877) );
  INV U6149 ( .IN(n5876), .OUT(n2685) );
  INV U6150 ( .IN(n5878), .OUT(n2688) );
  INV U6151 ( .IN(n4033), .OUT(n5880) );
  INV U6152 ( .IN(n5879), .OUT(n2691) );
  INV U6153 ( .IN(n5881), .OUT(n2694) );
  INV U6154 ( .IN(n4037), .OUT(n5883) );
  INV U6155 ( .IN(n5882), .OUT(n2697) );
  INV U6156 ( .IN(n5884), .OUT(n2700) );
  INV U6157 ( .IN(n4041), .OUT(n5886) );
  INV U6158 ( .IN(n5885), .OUT(n2703) );
  INV U6159 ( .IN(n6333), .OUT(n3456) );
  INV U6160 ( .IN(n4563), .OUT(n6362) );
  INV U6161 ( .IN(n6361), .OUT(n3459) );
  INV U6162 ( .IN(\mult_49/ab[1][20] ), .OUT(n1055) );
  INV U6163 ( .IN(n5888), .OUT(n2708) );
  INV U6164 ( .IN(n2707), .OUT(n5889) );
  INV U6165 ( .IN(n5891), .OUT(n2715) );
  INV U6166 ( .IN(n4050), .OUT(n5893) );
  INV U6167 ( .IN(n5892), .OUT(n2718) );
  INV U6168 ( .IN(n5894), .OUT(n2721) );
  INV U6169 ( .IN(n4054), .OUT(n5896) );
  INV U6170 ( .IN(n5895), .OUT(n2724) );
  INV U6171 ( .IN(n5897), .OUT(n2727) );
  INV U6172 ( .IN(n4058), .OUT(n5899) );
  INV U6173 ( .IN(n5898), .OUT(n2730) );
  INV U6174 ( .IN(n5900), .OUT(n2733) );
  INV U6175 ( .IN(n4062), .OUT(n5902) );
  INV U6176 ( .IN(n5901), .OUT(n2736) );
  INV U6177 ( .IN(n5903), .OUT(n2739) );
  INV U6178 ( .IN(n4066), .OUT(n5905) );
  INV U6179 ( .IN(n5904), .OUT(n2742) );
  INV U6180 ( .IN(n5906), .OUT(n2745) );
  INV U6181 ( .IN(n4070), .OUT(n5908) );
  INV U6182 ( .IN(n5907), .OUT(n2748) );
  INV U6183 ( .IN(n5909), .OUT(n2751) );
  INV U6184 ( .IN(n4074), .OUT(n5911) );
  INV U6185 ( .IN(n5910), .OUT(n2754) );
  INV U6186 ( .IN(n5912), .OUT(n2757) );
  INV U6187 ( .IN(n4526), .OUT(n6335) );
  INV U6188 ( .IN(n6334), .OUT(n3462) );
  INV U6189 ( .IN(n6363), .OUT(n3464) );
  INV U6190 ( .IN(\mult_49/ab[1][21] ), .OUT(n1131) );
  INV U6191 ( .IN(n5914), .OUT(n2762) );
  INV U6192 ( .IN(n2761), .OUT(n5915) );
  INV U6193 ( .IN(n5917), .OUT(n2769) );
  INV U6194 ( .IN(n4085), .OUT(n5919) );
  INV U6195 ( .IN(n5918), .OUT(n2772) );
  INV U6196 ( .IN(n5920), .OUT(n2775) );
  INV U6197 ( .IN(n4089), .OUT(n5922) );
  INV U6198 ( .IN(n5921), .OUT(n2778) );
  INV U6199 ( .IN(n5923), .OUT(n2781) );
  INV U6200 ( .IN(n4093), .OUT(n5925) );
  INV U6201 ( .IN(n5924), .OUT(n2784) );
  INV U6202 ( .IN(n5926), .OUT(n2787) );
  INV U6203 ( .IN(n4097), .OUT(n5928) );
  INV U6204 ( .IN(n5927), .OUT(n2790) );
  INV U6205 ( .IN(n5929), .OUT(n2793) );
  INV U6206 ( .IN(n4101), .OUT(n5931) );
  INV U6207 ( .IN(n5930), .OUT(n2796) );
  INV U6208 ( .IN(n5932), .OUT(n2799) );
  INV U6209 ( .IN(n4105), .OUT(n5934) );
  INV U6210 ( .IN(n5933), .OUT(n2802) );
  INV U6211 ( .IN(n5935), .OUT(n2805) );
  INV U6212 ( .IN(n4109), .OUT(n5937) );
  INV U6213 ( .IN(n5936), .OUT(n2808) );
  INV U6214 ( .IN(n5938), .OUT(n2811) );
  INV U6215 ( .IN(n4113), .OUT(n5940) );
  INV U6216 ( .IN(n5939), .OUT(n2814) );
  INV U6217 ( .IN(n6336), .OUT(n3468) );
  INV U6218 ( .IN(n4567), .OUT(n6365) );
  INV U6219 ( .IN(n6364), .OUT(n3471) );
  INV U6220 ( .IN(\mult_49/ab[1][22] ), .OUT(n1211) );
  INV U6221 ( .IN(n5942), .OUT(n2819) );
  INV U6222 ( .IN(n2818), .OUT(n5943) );
  INV U6223 ( .IN(n5945), .OUT(n2826) );
  INV U6224 ( .IN(n4122), .OUT(n5947) );
  INV U6225 ( .IN(n5946), .OUT(n2829) );
  INV U6226 ( .IN(n5948), .OUT(n2832) );
  INV U6227 ( .IN(n4126), .OUT(n5950) );
  INV U6228 ( .IN(n5949), .OUT(n2835) );
  INV U6229 ( .IN(n5951), .OUT(n2838) );
  INV U6230 ( .IN(n4130), .OUT(n5953) );
  INV U6231 ( .IN(n5952), .OUT(n2841) );
  INV U6232 ( .IN(n5954), .OUT(n2844) );
  INV U6233 ( .IN(n4134), .OUT(n5956) );
  INV U6234 ( .IN(n5955), .OUT(n2847) );
  INV U6235 ( .IN(n5957), .OUT(n2850) );
  INV U6236 ( .IN(n4138), .OUT(n5959) );
  INV U6237 ( .IN(n5958), .OUT(n2853) );
  INV U6238 ( .IN(n5960), .OUT(n2856) );
  INV U6239 ( .IN(n4142), .OUT(n5962) );
  INV U6240 ( .IN(n5961), .OUT(n2859) );
  INV U6241 ( .IN(n5963), .OUT(n2862) );
  INV U6242 ( .IN(n4146), .OUT(n5965) );
  INV U6243 ( .IN(n5964), .OUT(n2865) );
  INV U6244 ( .IN(n5966), .OUT(n2868) );
  INV U6245 ( .IN(n4150), .OUT(n5968) );
  INV U6246 ( .IN(n5967), .OUT(n2871) );
  INV U6247 ( .IN(n5969), .OUT(n2874) );
  INV U6248 ( .IN(n4530), .OUT(n6338) );
  INV U6249 ( .IN(n6337), .OUT(n3474) );
  INV U6250 ( .IN(n6366), .OUT(n3476) );
  INV U6251 ( .IN(\mult_49/ab[1][23] ), .OUT(n1295) );
  INV U6252 ( .IN(n5971), .OUT(n2879) );
  INV U6253 ( .IN(n2878), .OUT(n5972) );
  INV U6254 ( .IN(n5974), .OUT(n2886) );
  INV U6255 ( .IN(n4161), .OUT(n5976) );
  INV U6256 ( .IN(n5975), .OUT(n2889) );
  INV U6257 ( .IN(n5977), .OUT(n2892) );
  INV U6258 ( .IN(n4165), .OUT(n5979) );
  INV U6259 ( .IN(n5978), .OUT(n2895) );
  INV U6260 ( .IN(n5980), .OUT(n2898) );
  INV U6261 ( .IN(n4169), .OUT(n5982) );
  INV U6262 ( .IN(n5981), .OUT(n2901) );
  INV U6263 ( .IN(n5983), .OUT(n2904) );
  INV U6264 ( .IN(n4173), .OUT(n5985) );
  INV U6265 ( .IN(n5984), .OUT(n2907) );
  INV U6266 ( .IN(n5986), .OUT(n2910) );
  INV U6267 ( .IN(n4177), .OUT(n5988) );
  INV U6268 ( .IN(n5987), .OUT(n2913) );
  INV U6269 ( .IN(n5989), .OUT(n2916) );
  INV U6270 ( .IN(n4181), .OUT(n5991) );
  INV U6271 ( .IN(n5990), .OUT(n2919) );
  INV U6272 ( .IN(n5992), .OUT(n2922) );
  INV U6273 ( .IN(n4185), .OUT(n5994) );
  INV U6274 ( .IN(n5993), .OUT(n2925) );
  INV U6275 ( .IN(n5995), .OUT(n2928) );
  INV U6276 ( .IN(n4189), .OUT(n5997) );
  INV U6277 ( .IN(n5996), .OUT(n2931) );
  INV U6278 ( .IN(n5998), .OUT(n2934) );
  INV U6279 ( .IN(n4193), .OUT(n6000) );
  INV U6280 ( .IN(n5999), .OUT(n2937) );
  INV U6281 ( .IN(n6339), .OUT(n3480) );
  INV U6282 ( .IN(n4571), .OUT(n6368) );
  INV U6283 ( .IN(n6367), .OUT(n3483) );
  INV U6284 ( .IN(\mult_49/ab[1][24] ), .OUT(n1383) );
  INV U6285 ( .IN(n6002), .OUT(n2942) );
  INV U6286 ( .IN(n2941), .OUT(n6003) );
  INV U6287 ( .IN(n6005), .OUT(n2949) );
  INV U6288 ( .IN(n4202), .OUT(n6007) );
  INV U6289 ( .IN(n6006), .OUT(n2952) );
  INV U6290 ( .IN(n6008), .OUT(n2955) );
  INV U6291 ( .IN(n4206), .OUT(n6010) );
  INV U6292 ( .IN(n6009), .OUT(n2958) );
  INV U6293 ( .IN(n6011), .OUT(n2961) );
  INV U6294 ( .IN(n4210), .OUT(n6013) );
  INV U6295 ( .IN(n6012), .OUT(n2964) );
  INV U6296 ( .IN(n6014), .OUT(n2967) );
  INV U6297 ( .IN(n4214), .OUT(n6016) );
  INV U6298 ( .IN(n6015), .OUT(n2970) );
  INV U6299 ( .IN(n6017), .OUT(n2973) );
  INV U6300 ( .IN(n4218), .OUT(n6019) );
  INV U6301 ( .IN(n6018), .OUT(n2976) );
  INV U6302 ( .IN(n6020), .OUT(n2979) );
  INV U6303 ( .IN(n4222), .OUT(n6022) );
  INV U6304 ( .IN(n6021), .OUT(n2982) );
  INV U6305 ( .IN(n6023), .OUT(n2985) );
  INV U6306 ( .IN(n4226), .OUT(n6025) );
  INV U6307 ( .IN(n6024), .OUT(n2988) );
  INV U6308 ( .IN(n6026), .OUT(n2991) );
  INV U6309 ( .IN(n4230), .OUT(n6028) );
  INV U6310 ( .IN(n6027), .OUT(n2994) );
  INV U6311 ( .IN(n6029), .OUT(n2997) );
  INV U6312 ( .IN(n4234), .OUT(n6031) );
  INV U6313 ( .IN(n6030), .OUT(n3000) );
  INV U6314 ( .IN(n6032), .OUT(n3003) );
  INV U6315 ( .IN(n4534), .OUT(n6341) );
  INV U6316 ( .IN(n6340), .OUT(n3486) );
  INV U6317 ( .IN(n6369), .OUT(n3488) );
  INV U6318 ( .IN(\mult_49/ab[1][25] ), .OUT(n1475) );
  INV U6319 ( .IN(n6034), .OUT(n3008) );
  INV U6320 ( .IN(n3007), .OUT(n6035) );
  INV U6321 ( .IN(n6037), .OUT(n3015) );
  INV U6322 ( .IN(n4245), .OUT(n6039) );
  INV U6323 ( .IN(n6038), .OUT(n3018) );
  INV U6324 ( .IN(n6040), .OUT(n3021) );
  INV U6325 ( .IN(n4249), .OUT(n6042) );
  INV U6326 ( .IN(n6041), .OUT(n3024) );
  INV U6327 ( .IN(n6043), .OUT(n3027) );
  INV U6328 ( .IN(n4253), .OUT(n6045) );
  INV U6329 ( .IN(n6044), .OUT(n3030) );
  INV U6330 ( .IN(n6046), .OUT(n3033) );
  INV U6331 ( .IN(n4257), .OUT(n6048) );
  INV U6332 ( .IN(n6047), .OUT(n3036) );
  INV U6333 ( .IN(n6049), .OUT(n3039) );
  INV U6334 ( .IN(n4261), .OUT(n6051) );
  INV U6335 ( .IN(n6050), .OUT(n3042) );
  INV U6336 ( .IN(n6052), .OUT(n3045) );
  INV U6337 ( .IN(n4265), .OUT(n6054) );
  INV U6338 ( .IN(n6053), .OUT(n3048) );
  INV U6339 ( .IN(n6055), .OUT(n3051) );
  INV U6340 ( .IN(n4269), .OUT(n6057) );
  INV U6341 ( .IN(n6056), .OUT(n3054) );
  INV U6342 ( .IN(n6058), .OUT(n3057) );
  INV U6343 ( .IN(n4273), .OUT(n6060) );
  INV U6344 ( .IN(n6059), .OUT(n3060) );
  INV U6345 ( .IN(n6061), .OUT(n3063) );
  INV U6346 ( .IN(n4277), .OUT(n6063) );
  INV U6347 ( .IN(n6062), .OUT(n3066) );
  INV U6348 ( .IN(n6064), .OUT(n3069) );
  INV U6349 ( .IN(n4281), .OUT(n6066) );
  INV U6350 ( .IN(n6065), .OUT(n3072) );
  INV U6351 ( .IN(n6342), .OUT(n3492) );
  INV U6352 ( .IN(n4575), .OUT(n6371) );
  INV U6353 ( .IN(n6370), .OUT(n3495) );
  INV U6354 ( .IN(\mult_49/ab[1][26] ), .OUT(n1571) );
  INV U6355 ( .IN(n6068), .OUT(n3077) );
  INV U6356 ( .IN(n3076), .OUT(n6069) );
  INV U6357 ( .IN(n6071), .OUT(n3084) );
  INV U6358 ( .IN(n4290), .OUT(n6073) );
  INV U6359 ( .IN(n6072), .OUT(n3087) );
  INV U6360 ( .IN(n6074), .OUT(n3090) );
  INV U6361 ( .IN(n4294), .OUT(n6076) );
  INV U6362 ( .IN(n6075), .OUT(n3093) );
  INV U6363 ( .IN(n6077), .OUT(n3096) );
  INV U6364 ( .IN(n4298), .OUT(n6079) );
  INV U6365 ( .IN(n6078), .OUT(n3099) );
  INV U6366 ( .IN(n6080), .OUT(n3102) );
  INV U6367 ( .IN(n4302), .OUT(n6082) );
  INV U6368 ( .IN(n6081), .OUT(n3105) );
  INV U6369 ( .IN(n6083), .OUT(n3108) );
  INV U6370 ( .IN(n4306), .OUT(n6085) );
  INV U6371 ( .IN(n6084), .OUT(n3111) );
  INV U6372 ( .IN(n6086), .OUT(n3114) );
  INV U6373 ( .IN(n4310), .OUT(n6088) );
  INV U6374 ( .IN(n6087), .OUT(n3117) );
  INV U6375 ( .IN(n6089), .OUT(n3120) );
  INV U6376 ( .IN(n4314), .OUT(n6091) );
  INV U6377 ( .IN(n6090), .OUT(n3123) );
  INV U6378 ( .IN(n6092), .OUT(n3126) );
  INV U6379 ( .IN(n4318), .OUT(n6094) );
  INV U6380 ( .IN(n6093), .OUT(n3129) );
  INV U6381 ( .IN(n6095), .OUT(n3132) );
  INV U6382 ( .IN(n4322), .OUT(n6097) );
  INV U6383 ( .IN(n6096), .OUT(n3135) );
  INV U6384 ( .IN(n6098), .OUT(n3138) );
  INV U6385 ( .IN(n4326), .OUT(n6100) );
  INV U6386 ( .IN(n6099), .OUT(n3141) );
  INV U6387 ( .IN(n6101), .OUT(n3144) );
  INV U6388 ( .IN(n4538), .OUT(n6344) );
  INV U6389 ( .IN(n6343), .OUT(n3498) );
  INV U6390 ( .IN(n6372), .OUT(n3500) );
  INV U6391 ( .IN(\mult_49/ab[1][27] ), .OUT(n1671) );
  INV U6392 ( .IN(n6103), .OUT(n3149) );
  INV U6393 ( .IN(n3148), .OUT(n6104) );
  INV U6394 ( .IN(n6106), .OUT(n3156) );
  INV U6395 ( .IN(n4337), .OUT(n6108) );
  INV U6396 ( .IN(n6107), .OUT(n3159) );
  INV U6397 ( .IN(n6109), .OUT(n3162) );
  INV U6398 ( .IN(n4341), .OUT(n6111) );
  INV U6399 ( .IN(n6110), .OUT(n3165) );
  INV U6400 ( .IN(n6112), .OUT(n3168) );
  INV U6401 ( .IN(n4345), .OUT(n6114) );
  INV U6402 ( .IN(n6113), .OUT(n3171) );
  INV U6403 ( .IN(n6115), .OUT(n3174) );
  INV U6404 ( .IN(n4349), .OUT(n6117) );
  INV U6405 ( .IN(n6116), .OUT(n3177) );
  INV U6406 ( .IN(n6118), .OUT(n3180) );
  INV U6407 ( .IN(n4353), .OUT(n6120) );
  INV U6408 ( .IN(n6119), .OUT(n3183) );
  INV U6409 ( .IN(n6121), .OUT(n3186) );
  INV U6410 ( .IN(n4357), .OUT(n6123) );
  INV U6411 ( .IN(n6122), .OUT(n3189) );
  INV U6412 ( .IN(n6124), .OUT(n3192) );
  INV U6413 ( .IN(n4361), .OUT(n6126) );
  INV U6414 ( .IN(n6125), .OUT(n3195) );
  INV U6415 ( .IN(n6127), .OUT(n3198) );
  INV U6416 ( .IN(n4365), .OUT(n6129) );
  INV U6417 ( .IN(n6128), .OUT(n3201) );
  INV U6418 ( .IN(n6130), .OUT(n3204) );
  INV U6419 ( .IN(n4369), .OUT(n6132) );
  INV U6420 ( .IN(n6131), .OUT(n3207) );
  INV U6421 ( .IN(n6133), .OUT(n3210) );
  INV U6422 ( .IN(n4373), .OUT(n6135) );
  INV U6423 ( .IN(n6134), .OUT(n3213) );
  INV U6424 ( .IN(n6136), .OUT(n3216) );
  INV U6425 ( .IN(n4377), .OUT(n6138) );
  INV U6426 ( .IN(n6137), .OUT(n3219) );
  INV U6427 ( .IN(n6345), .OUT(n3504) );
  INV U6428 ( .IN(n4579), .OUT(n6374) );
  INV U6429 ( .IN(n6373), .OUT(n3507) );
  INV U6430 ( .IN(\mult_49/ab[1][28] ), .OUT(n1775) );
  INV U6431 ( .IN(n6140), .OUT(n3224) );
  INV U6432 ( .IN(n3223), .OUT(n6141) );
  INV U6433 ( .IN(n6143), .OUT(n3231) );
  INV U6434 ( .IN(n4386), .OUT(n6145) );
  INV U6435 ( .IN(n6144), .OUT(n3234) );
  INV U6436 ( .IN(n6146), .OUT(n3237) );
  INV U6437 ( .IN(n4390), .OUT(n6148) );
  INV U6438 ( .IN(n6147), .OUT(n3240) );
  INV U6439 ( .IN(n6149), .OUT(n3243) );
  INV U6440 ( .IN(n4394), .OUT(n6151) );
  INV U6441 ( .IN(n6150), .OUT(n3246) );
  INV U6442 ( .IN(n6152), .OUT(n3249) );
  INV U6443 ( .IN(n4398), .OUT(n6154) );
  INV U6444 ( .IN(n6153), .OUT(n3252) );
  INV U6445 ( .IN(n6155), .OUT(n3255) );
  INV U6446 ( .IN(n4402), .OUT(n6157) );
  INV U6447 ( .IN(n6156), .OUT(n3258) );
  INV U6448 ( .IN(n6158), .OUT(n3261) );
  INV U6449 ( .IN(n4406), .OUT(n6160) );
  INV U6450 ( .IN(n6159), .OUT(n3264) );
  INV U6451 ( .IN(n6161), .OUT(n3267) );
  INV U6452 ( .IN(n4410), .OUT(n6163) );
  INV U6453 ( .IN(n6162), .OUT(n3270) );
  INV U6454 ( .IN(n6164), .OUT(n3273) );
  INV U6455 ( .IN(n4414), .OUT(n6166) );
  INV U6456 ( .IN(n6165), .OUT(n3276) );
  INV U6457 ( .IN(n6167), .OUT(n3279) );
  INV U6458 ( .IN(n4418), .OUT(n6169) );
  INV U6459 ( .IN(n6168), .OUT(n3282) );
  INV U6460 ( .IN(n6170), .OUT(n3285) );
  INV U6461 ( .IN(n4422), .OUT(n6172) );
  INV U6462 ( .IN(n6171), .OUT(n3288) );
  INV U6463 ( .IN(n6173), .OUT(n3291) );
  INV U6464 ( .IN(n4426), .OUT(n6175) );
  INV U6465 ( .IN(n6174), .OUT(n3294) );
  INV U6466 ( .IN(n6176), .OUT(n3297) );
  INV U6467 ( .IN(n4542), .OUT(n6347) );
  INV U6468 ( .IN(n6346), .OUT(n3510) );
  INV U6469 ( .IN(n6375), .OUT(n3512) );
  INV U6470 ( .IN(n6177), .OUT(n3300) );
  INV U6471 ( .IN(n6179), .OUT(n3303) );
  INV U6472 ( .IN(n3301), .OUT(n6180) );
  INV U6473 ( .IN(n6182), .OUT(n3309) );
  INV U6474 ( .IN(n4439), .OUT(n6184) );
  INV U6475 ( .IN(n6183), .OUT(n3312) );
  INV U6476 ( .IN(n6185), .OUT(n3315) );
  INV U6477 ( .IN(n4445), .OUT(n6187) );
  INV U6478 ( .IN(n6186), .OUT(n3318) );
  INV U6479 ( .IN(n6188), .OUT(n3321) );
  INV U6480 ( .IN(n4451), .OUT(n6190) );
  INV U6481 ( .IN(n6189), .OUT(n3324) );
  INV U6482 ( .IN(n6191), .OUT(n3327) );
  INV U6483 ( .IN(n4457), .OUT(n6193) );
  INV U6484 ( .IN(n6192), .OUT(n3330) );
  INV U6485 ( .IN(n6194), .OUT(n3333) );
  INV U6486 ( .IN(n4463), .OUT(n6196) );
  INV U6487 ( .IN(n6195), .OUT(n3336) );
  INV U6488 ( .IN(n6197), .OUT(n3339) );
  INV U6489 ( .IN(n4469), .OUT(n6199) );
  INV U6490 ( .IN(n6198), .OUT(n3342) );
  INV U6491 ( .IN(n6200), .OUT(n3345) );
  INV U6492 ( .IN(n4475), .OUT(n6202) );
  INV U6493 ( .IN(n6201), .OUT(n3348) );
  INV U6494 ( .IN(n6203), .OUT(n3351) );
  INV U6495 ( .IN(n4481), .OUT(n6205) );
  INV U6496 ( .IN(n6204), .OUT(n3354) );
  INV U6497 ( .IN(n6206), .OUT(n3357) );
  INV U6498 ( .IN(n4487), .OUT(n6208) );
  INV U6499 ( .IN(n6207), .OUT(n3360) );
  INV U6500 ( .IN(n6209), .OUT(n3363) );
  INV U6501 ( .IN(n4493), .OUT(n6211) );
  INV U6502 ( .IN(n6210), .OUT(n3366) );
  INV U6503 ( .IN(n6212), .OUT(n3369) );
  INV U6504 ( .IN(n4499), .OUT(n6214) );
  INV U6505 ( .IN(n6213), .OUT(n3372) );
  INV U6506 ( .IN(n6215), .OUT(n3375) );
  INV U6507 ( .IN(n4505), .OUT(n6217) );
  INV U6508 ( .IN(n6216), .OUT(n3378) );
  INV U6509 ( .IN(n6348), .OUT(n3516) );
  INV U6510 ( .IN(n4583), .OUT(n6377) );
  INV U6511 ( .IN(n6376), .OUT(n3519) );
  INV U6512 ( .IN(n6378), .OUT(n4723) );
  INV U6513 ( .IN(n6316), .OUT(n4708) );
  INV U6514 ( .IN(n6310), .OUT(n4678) );
  INV U6515 ( .IN(n6307), .OUT(n4675) );
  INV U6516 ( .IN(n6311), .OUT(n3399) );
  INV U6517 ( .IN(n6302), .OUT(n4669) );
  INV U6518 ( .IN(n6296), .OUT(n4639) );
  INV U6519 ( .IN(n6293), .OUT(n4636) );
  INV U6520 ( .IN(n6297), .OUT(n3390) );
  INV U6521 ( .IN(n6288), .OUT(n4630) );
  INV U6522 ( .IN(n6283), .OUT(n4615) );
  INV U6523 ( .IN(n6278), .OUT(n4600) );
  INV U6524 ( .IN(n6275), .OUT(n4597) );
  INV U6525 ( .IN(n6280), .OUT(n4603) );
  INV U6526 ( .IN(n6272), .OUT(n4590) );
  INV U6527 ( .IN(n6269), .OUT(n4588) );
  INV U6528 ( .IN(n6273), .OUT(n4594) );
  INV U6529 ( .IN(n6281), .OUT(n3381) );
  INV U6530 ( .IN(n6285), .OUT(n4618) );
  INV U6531 ( .IN(n6266), .OUT(n4609) );
  INV U6532 ( .IN(n6263), .OUT(n4606) );
  INV U6533 ( .IN(n6267), .OUT(n4612) );
  INV U6534 ( .IN(n6286), .OUT(n3384) );
  INV U6535 ( .IN(n6290), .OUT(n4633) );
  INV U6536 ( .IN(n6259), .OUT(n4624) );
  INV U6537 ( .IN(n6256), .OUT(n4621) );
  INV U6538 ( .IN(n6261), .OUT(n4627) );
  INV U6539 ( .IN(n6291), .OUT(n3387) );
  INV U6540 ( .IN(n6298), .OUT(n4654) );
  INV U6541 ( .IN(n6253), .OUT(n4651) );
  INV U6542 ( .IN(n6299), .OUT(n4657) );
  INV U6543 ( .IN(n6250), .OUT(n4645) );
  INV U6544 ( .IN(n6247), .OUT(n4642) );
  INV U6545 ( .IN(n6251), .OUT(n4648) );
  INV U6546 ( .IN(n6300), .OUT(n3393) );
  INV U6547 ( .IN(n6304), .OUT(n4672) );
  INV U6548 ( .IN(n6243), .OUT(n4663) );
  INV U6549 ( .IN(n6240), .OUT(n4660) );
  INV U6550 ( .IN(n6245), .OUT(n4666) );
  INV U6551 ( .IN(n6305), .OUT(n3396) );
  INV U6552 ( .IN(n6312), .OUT(n4693) );
  INV U6553 ( .IN(n6237), .OUT(n4690) );
  INV U6554 ( .IN(n6313), .OUT(n4696) );
  INV U6555 ( .IN(n6234), .OUT(n4684) );
  INV U6556 ( .IN(n6231), .OUT(n4681) );
  INV U6557 ( .IN(n6235), .OUT(n4687) );
  INV U6558 ( .IN(n6314), .OUT(n3402) );
  INV U6559 ( .IN(n6318), .OUT(n4711) );
  INV U6560 ( .IN(n6227), .OUT(n4702) );
  INV U6561 ( .IN(n6224), .OUT(n4699) );
  INV U6562 ( .IN(n6229), .OUT(n4705) );
  INV U6563 ( .IN(n6319), .OUT(n3405) );
  INV U6564 ( .IN(n6380), .OUT(n4726) );
  INV U6565 ( .IN(n6221), .OUT(n4717) );
  INV U6566 ( .IN(n6218), .OUT(n4714) );
  INV U6567 ( .IN(n6222), .OUT(n4720) );
  INV U6568 ( .IN(n6381), .OUT(n3521) );
  INV U6569 ( .IN(\mult_49/ab[29][2] ), .OUT(n5715) );
  INV U6570 ( .IN(n4856), .OUT(n4857) );
  INV U6571 ( .IN(n4859), .OUT(n4860) );
  INV U6572 ( .IN(n4862), .OUT(n4863) );
  INV U6573 ( .IN(n4865), .OUT(n4866) );
  INV U6574 ( .IN(n4755), .OUT(n4870) );
  INV U6575 ( .IN(n4872), .OUT(n4873) );
  INV U6576 ( .IN(n4875), .OUT(n4876) );
  INV U6577 ( .IN(n4878), .OUT(n4879) );
  INV U6578 ( .IN(n4881), .OUT(n4882) );
  INV U6579 ( .IN(n4884), .OUT(n4885) );
  INV U6580 ( .IN(n6394), .OUT(n3543) );
  INV U6581 ( .IN(n6395), .OUT(n3567) );
  INV U6582 ( .IN(n4890), .OUT(n4891) );
  INV U6583 ( .IN(n4896), .OUT(n4897) );
  INV U6584 ( .IN(n4902), .OUT(n4903) );
  INV U6585 ( .IN(n4908), .OUT(n4909) );
  INV U6586 ( .IN(n4914), .OUT(n4915) );
  INV U6587 ( .IN(n2091), .OUT(n6397) );
  INV U6588 ( .IN(n6398), .OUT(n3642) );
  INV U6589 ( .IN(n4924), .OUT(n4925) );
  INV U6590 ( .IN(n4930), .OUT(n4931) );
  INV U6591 ( .IN(n4936), .OUT(n4937) );
  INV U6592 ( .IN(n4942), .OUT(n4943) );
  INV U6593 ( .IN(n4948), .OUT(n4949) );
  INV U6594 ( .IN(n4954), .OUT(n4955) );
  INV U6595 ( .IN(n4960), .OUT(n4961) );
  INV U6596 ( .IN(n4966), .OUT(n4967) );
  INV U6597 ( .IN(n4972), .OUT(n4973) );
  INV U6598 ( .IN(n4978), .OUT(n4979) );
  INV U6599 ( .IN(n4984), .OUT(n4985) );
  INV U6600 ( .IN(n4990), .OUT(n4991) );
  INV U6601 ( .IN(n4996), .OUT(n4997) );
  INV U6602 ( .IN(n5002), .OUT(n5003) );
  INV U6603 ( .IN(n5008), .OUT(n5009) );
  INV U6604 ( .IN(n5014), .OUT(n5015) );
  INV U6605 ( .IN(n5020), .OUT(n5021) );
  INV U6606 ( .IN(n5026), .OUT(n5027) );
  INV U6607 ( .IN(n5032), .OUT(n5033) );
  INV U6608 ( .IN(n5038), .OUT(n5039) );
  INV U6609 ( .IN(n5044), .OUT(n5045) );
  INV U6610 ( .IN(n5050), .OUT(n5051) );
  INV U6611 ( .IN(n5056), .OUT(n5057) );
  INV U6612 ( .IN(n5062), .OUT(n5063) );
  INV U6613 ( .IN(n5068), .OUT(n5069) );
  INV U6614 ( .IN(n6399), .OUT(\gt_48/LTV1 [31]) );
  INV U6615 ( .IN(\gt_48/SB ), .OUT(n6400) );
  INV U6616 ( .IN(n6401), .OUT(\gt_48/LTV1 [30]) );
  INV U6617 ( .IN(A[30]), .OUT(n6402) );
  INV U6618 ( .IN(n6403), .OUT(\gt_48/LTV1 [29]) );
  INV U6619 ( .IN(A[29]), .OUT(n6404) );
  INV U6620 ( .IN(n6405), .OUT(\gt_48/LTV1 [28]) );
  INV U6621 ( .IN(A[28]), .OUT(n6406) );
  INV U6622 ( .IN(n6407), .OUT(\gt_48/LTV1 [27]) );
  INV U6623 ( .IN(A[27]), .OUT(n6408) );
  INV U6624 ( .IN(n6409), .OUT(\gt_48/LTV1 [26]) );
  INV U6625 ( .IN(A[26]), .OUT(n6410) );
  INV U6626 ( .IN(n6411), .OUT(\gt_48/LTV1 [25]) );
  INV U6627 ( .IN(A[25]), .OUT(n6412) );
  INV U6628 ( .IN(n6413), .OUT(\gt_48/LTV1 [24]) );
  INV U6629 ( .IN(A[24]), .OUT(n6414) );
  INV U6630 ( .IN(n6415), .OUT(\gt_48/LTV1 [23]) );
  INV U6631 ( .IN(A[23]), .OUT(n6416) );
  INV U6632 ( .IN(n6417), .OUT(\gt_48/LTV1 [22]) );
  INV U6633 ( .IN(A[22]), .OUT(n6418) );
  INV U6634 ( .IN(n6419), .OUT(\gt_48/LTV1 [21]) );
  INV U6635 ( .IN(A[21]), .OUT(n6420) );
  INV U6636 ( .IN(n6421), .OUT(\gt_48/LTV1 [20]) );
  INV U6637 ( .IN(A[20]), .OUT(n6422) );
  INV U6638 ( .IN(n6423), .OUT(\gt_48/LTV1 [19]) );
  INV U6639 ( .IN(A[19]), .OUT(n6424) );
  INV U6640 ( .IN(n6425), .OUT(\gt_48/LTV1 [18]) );
  INV U6641 ( .IN(A[18]), .OUT(n6426) );
  INV U6642 ( .IN(n6427), .OUT(\gt_48/LTV1 [17]) );
  INV U6643 ( .IN(A[17]), .OUT(n6428) );
  INV U6644 ( .IN(n6429), .OUT(\gt_48/LTV1 [16]) );
  INV U6645 ( .IN(A[16]), .OUT(n6430) );
  INV U6646 ( .IN(n6431), .OUT(\gt_48/LTV1 [15]) );
  INV U6647 ( .IN(A[15]), .OUT(n6432) );
  INV U6648 ( .IN(n6433), .OUT(\gt_48/LTV1 [14]) );
  INV U6649 ( .IN(A[14]), .OUT(n6434) );
  INV U6650 ( .IN(n6435), .OUT(\gt_48/LTV1 [13]) );
  INV U6651 ( .IN(A[13]), .OUT(n6436) );
  INV U6652 ( .IN(n6437), .OUT(\gt_48/LTV1 [12]) );
  INV U6653 ( .IN(A[12]), .OUT(n6438) );
  INV U6654 ( .IN(n6439), .OUT(\gt_48/LTV1 [11]) );
  INV U6655 ( .IN(A[11]), .OUT(n6440) );
  INV U6656 ( .IN(n6441), .OUT(\gt_48/LTV1 [10]) );
  INV U6657 ( .IN(A[10]), .OUT(n6442) );
  INV U6658 ( .IN(n6443), .OUT(\gt_48/LTV1 [9]) );
  INV U6659 ( .IN(A[9]), .OUT(n6444) );
  INV U6660 ( .IN(n6445), .OUT(\gt_48/LTV1 [8]) );
  INV U6661 ( .IN(A[8]), .OUT(n6446) );
  INV U6662 ( .IN(n6447), .OUT(\gt_48/LTV1 [7]) );
  INV U6663 ( .IN(A[7]), .OUT(n6448) );
  INV U6664 ( .IN(n6449), .OUT(\gt_48/LTV1 [6]) );
  INV U6665 ( .IN(A[6]), .OUT(n6450) );
  INV U6666 ( .IN(n6451), .OUT(\gt_48/LTV1 [5]) );
  INV U6667 ( .IN(A[5]), .OUT(n6452) );
  INV U6668 ( .IN(n6453), .OUT(\gt_48/LTV1 [4]) );
  INV U6669 ( .IN(A[4]), .OUT(n6454) );
  INV U6670 ( .IN(n6455), .OUT(\gt_48/LTV1 [3]) );
  INV U6671 ( .IN(A[3]), .OUT(n6456) );
  INV U6672 ( .IN(n6457), .OUT(\gt_48/LTV1 [2]) );
  INV U6673 ( .IN(A[2]), .OUT(n6458) );
  INV U6674 ( .IN(n6459), .OUT(\gt_48/LTV1 [1]) );
  INV U6675 ( .IN(A[1]), .OUT(n6460) );
  INV U6676 ( .IN(n6461), .OUT(\gt_48/LTV1 [0]) );
  INV U6677 ( .IN(A[0]), .OUT(n6462) );
endmodule

